/*
[Bare framework] Leave empty, this is used when exporting to verilog
*/

module M_mul_cmp16_0_M_frame_display_div_mc0 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>0);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_0_M_frame_display_div_mc1 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>0);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_0_M_frame_display_div_mc2 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>0);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_0_M_frame_display_div_mc3 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>0);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_0_M_frame_display_div_mc4 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>0);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_0_M_frame_display_div_mc5 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>0);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_0_M_frame_display_div_mc6 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>0);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_0_M_frame_display_div_mc7 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>0);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_8_M_frame_display_div_mc8 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>8);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_8_M_frame_display_div_mc9 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>8);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_8_M_frame_display_div_mc10 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>8);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_8_M_frame_display_div_mc11 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>8);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_8_M_frame_display_div_mc12 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>8);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_8_M_frame_display_div_mc13 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>8);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_mul_cmp16_8_M_frame_display_div_mc14 (
in_num,
in_den,
out_beq,
out_clock,
clock
);
input  [15:0] in_num;
input  [15:0] in_den;
output  [0:0] out_beq;
output out_clock;
input clock;
assign out_clock = clock;
reg  [16:0] _t_nk;
reg  [0:0] _t_beq;

assign out_beq = _t_beq;



`ifdef FORMAL
initial begin
assume(reset);
end
`endif
always @* begin
// _always_pre
// __block_1
_t_nk = (in_num>>8);

_t_beq = (_t_nk>in_den);

// __block_2
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
end

endmodule


module M_div16_M_frame_display_div (
in_inum,
in_iden,
out_ret,
in_run,
out_done,
reset,
out_clock,
clock
);
input signed [15:0] in_inum;
input signed [15:0] in_iden;
output signed [15:0] out_ret;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire  [0:0] _w_mc0_beq;
wire  [0:0] _w_mc1_beq;
wire  [0:0] _w_mc2_beq;
wire  [0:0] _w_mc3_beq;
wire  [0:0] _w_mc4_beq;
wire  [0:0] _w_mc5_beq;
wire  [0:0] _w_mc6_beq;
wire  [0:0] _w_mc7_beq;
wire  [0:0] _w_mc8_beq;
wire  [0:0] _w_mc9_beq;
wire  [0:0] _w_mc10_beq;
wire  [0:0] _w_mc11_beq;
wire  [0:0] _w_mc12_beq;
wire  [0:0] _w_mc13_beq;
wire  [0:0] _w_mc14_beq;
wire  [0:0] _c_num_neg;
assign _c_num_neg = 0;
wire  [0:0] _c_den_neg;
assign _c_den_neg = 0;
reg  [15:0] _t_num;
reg  [15:0] _t_concat;

reg  [15:0] _d_reminder;
reg  [15:0] _q_reminder;
reg  [15:0] _d_den;
reg  [15:0] _q_den;
reg signed [15:0] _d_ret;
reg signed [15:0] _q_ret;
reg  [1:0] _d__idx_fsm0,_q__idx_fsm0;
assign out_ret = _q_ret;
assign out_done = (_q__idx_fsm0 == 0)
;
M_mul_cmp16_0_M_frame_display_div_mc0 mc0 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc0_beq),
.clock(clock));
M_mul_cmp16_0_M_frame_display_div_mc1 mc1 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc1_beq),
.clock(clock));
M_mul_cmp16_0_M_frame_display_div_mc2 mc2 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc2_beq),
.clock(clock));
M_mul_cmp16_0_M_frame_display_div_mc3 mc3 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc3_beq),
.clock(clock));
M_mul_cmp16_0_M_frame_display_div_mc4 mc4 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc4_beq),
.clock(clock));
M_mul_cmp16_0_M_frame_display_div_mc5 mc5 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc5_beq),
.clock(clock));
M_mul_cmp16_0_M_frame_display_div_mc6 mc6 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc6_beq),
.clock(clock));
M_mul_cmp16_0_M_frame_display_div_mc7 mc7 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc7_beq),
.clock(clock));
M_mul_cmp16_8_M_frame_display_div_mc8 mc8 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc8_beq),
.clock(clock));
M_mul_cmp16_8_M_frame_display_div_mc9 mc9 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc9_beq),
.clock(clock));
M_mul_cmp16_8_M_frame_display_div_mc10 mc10 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc10_beq),
.clock(clock));
M_mul_cmp16_8_M_frame_display_div_mc11 mc11 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc11_beq),
.clock(clock));
M_mul_cmp16_8_M_frame_display_div_mc12 mc12 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc12_beq),
.clock(clock));
M_mul_cmp16_8_M_frame_display_div_mc13 mc13 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc13_beq),
.clock(clock));
M_mul_cmp16_8_M_frame_display_div_mc14 mc14 (
.in_num(_q_reminder),
.in_den(_q_den),
.out_beq(_w_mc14_beq),
.clock(clock));



`ifdef FORMAL
initial begin
assume(reset);
end
assume property($initstate || (in_run || out_done));
`endif
always @* begin
_d_reminder = _q_reminder;
_d_den = _q_den;
_d_ret = _q_ret;
_d__idx_fsm0 = _q__idx_fsm0;
_t_num = 0;
_t_concat = 0;
// _always_pre
(* full_case *)
case (_q__idx_fsm0)
1: begin
// _top
_d_den = in_iden;

_t_num = in_inum;

if (_d_den>_t_num) begin
// __block_1
// __block_3
_d_ret = 0;

_d__idx_fsm0 = 0;
end else begin
// __block_2
// collapsed 'after'
// __block_6
if (_d_den==_t_num) begin
// __block_7
// __block_9
_d_ret = 1;

_d__idx_fsm0 = 0;
end else begin
// __block_8
// collapsed 'after'
// __block_12
if (_d_den==0) begin
// __block_13
// __block_15
if (_c_num_neg^_c_den_neg) begin
// __block_16
// __block_18
_d_ret = 16'b1111111111111111;

// __block_19
end else begin
// __block_17
// __block_20
_d_ret = 16'b0111111111111111;

// __block_21
end
// 'after'
// __block_22
_d__idx_fsm0 = 0;
end else begin
// __block_14
// collapsed 'after'
// __block_25
_d_reminder = _t_num;

_d_ret = 0;

_d__idx_fsm0 = 3;
end
end
end
end
2: begin
// done
_d__idx_fsm0 = 0;
end
3: begin
// __while__block_26
if (_q_reminder>=_q_den) begin
// __block_27
// __block_29
_t_concat = {!_w_mc14_beq&&_w_mc13_beq,!_w_mc13_beq&&_w_mc12_beq,!_w_mc12_beq&&_w_mc11_beq,!_w_mc11_beq&&_w_mc10_beq,!_w_mc10_beq&&_w_mc9_beq,!_w_mc9_beq&&_w_mc8_beq,!_w_mc8_beq&&_w_mc7_beq,!_w_mc7_beq&&_w_mc6_beq,!_w_mc6_beq&&_w_mc5_beq,!_w_mc5_beq&&_w_mc4_beq,!_w_mc4_beq&&_w_mc3_beq,!_w_mc3_beq&&_w_mc2_beq,!_w_mc2_beq&&_w_mc1_beq,!_w_mc1_beq&&_w_mc0_beq,1'b0};

  case (_t_concat)
  16'b1000000000000000: begin
// __block_31_case
// __block_32
_d_ret = _q_ret+(1<<8);

_d_reminder = _q_reminder-(_q_den<<8);

// __block_33
  end
  16'b0100000000000000: begin
// __block_34_case
// __block_35
_d_ret = _q_ret+(1<<8);

_d_reminder = _q_reminder-(_q_den<<8);

// __block_36
  end
  16'b0010000000000000: begin
// __block_37_case
// __block_38
_d_ret = _q_ret+(1<<8);

_d_reminder = _q_reminder-(_q_den<<8);

// __block_39
  end
  16'b0001000000000000: begin
// __block_40_case
// __block_41
_d_ret = _q_ret+(1<<8);

_d_reminder = _q_reminder-(_q_den<<8);

// __block_42
  end
  16'b0000100000000000: begin
// __block_43_case
// __block_44
_d_ret = _q_ret+(1<<8);

_d_reminder = _q_reminder-(_q_den<<8);

// __block_45
  end
  16'b0000010000000000: begin
// __block_46_case
// __block_47
_d_ret = _q_ret+(1<<8);

_d_reminder = _q_reminder-(_q_den<<8);

// __block_48
  end
  16'b0000001000000000: begin
// __block_49_case
// __block_50
_d_ret = _q_ret+(1<<8);

_d_reminder = _q_reminder-(_q_den<<8);

// __block_51
  end
  16'b0000000100000000: begin
// __block_52_case
// __block_53
_d_ret = _q_ret+(1<<0);

_d_reminder = _q_reminder-(_q_den<<0);

// __block_54
  end
  16'b0000000010000000: begin
// __block_55_case
// __block_56
_d_ret = _q_ret+(1<<0);

_d_reminder = _q_reminder-(_q_den<<0);

// __block_57
  end
  16'b0000000001000000: begin
// __block_58_case
// __block_59
_d_ret = _q_ret+(1<<0);

_d_reminder = _q_reminder-(_q_den<<0);

// __block_60
  end
  16'b0000000000100000: begin
// __block_61_case
// __block_62
_d_ret = _q_ret+(1<<0);

_d_reminder = _q_reminder-(_q_den<<0);

// __block_63
  end
  16'b0000000000010000: begin
// __block_64_case
// __block_65
_d_ret = _q_ret+(1<<0);

_d_reminder = _q_reminder-(_q_den<<0);

// __block_66
  end
  16'b0000000000001000: begin
// __block_67_case
// __block_68
_d_ret = _q_ret+(1<<0);

_d_reminder = _q_reminder-(_q_den<<0);

// __block_69
  end
  16'b0000000000000100: begin
// __block_70_case
// __block_71
_d_ret = _q_ret+(1<<0);

_d_reminder = _q_reminder-(_q_den<<0);

// __block_72
  end
  16'b0000000000000010: begin
// __block_73_case
// __block_74
_d_ret = _q_ret+(1<<0);

_d_reminder = _q_reminder-(_q_den<<0);

// __block_75
  end
  16'b0000000000000000: begin
// __block_76_case
// __block_77
_d_ret = _q_ret+(1<<0);

_d_reminder = _q_reminder-(_q_den<<0);

// __block_78
  end
  default: begin
// __block_79_case
// __block_80
// __block_81
  end
endcase
// __block_30
// __block_82
_d__idx_fsm0 = 3;
end else begin
// __block_28
_d__idx_fsm0 = 0;
end
end
0: begin 
end
default: begin 
_d__idx_fsm0 = {2{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
_q_reminder <= (reset | ~in_run) ? 0 : _d_reminder;
_q_den <= (reset | ~in_run) ? 0 : _d_den;
_q_ret <= _d_ret;
_q__idx_fsm0 <= reset ? 0 : ( ~in_run ? 1 : _d__idx_fsm0);
end

endmodule


module M_frame_display (
in_pix_x,
in_pix_y,
in_pix_active,
in_pix_vblank,
in_vga_hs,
in_vga_vs,
out_pix_r,
out_pix_g,
out_pix_b,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [10:0] in_pix_x;
input  [10:0] in_pix_y;
input  [0:0] in_pix_active;
input  [0:0] in_pix_vblank;
input  [0:0] in_vga_hs;
input  [0:0] in_vga_vs;
output  [7:0] out_pix_r;
output  [7:0] out_pix_g;
output  [7:0] out_pix_b;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire signed [15:0] _w_div_ret;
wire _w_div_done;
wire  [14:0] _c_maxv;
assign _c_maxv = 22000;
reg  [8:0] _t_offs_y;
reg  [7:0] _t_u;
reg  [7:0] _t_v;
reg  [0:0] _t_floor;
reg  [7:0] _t_pix_r;
reg  [7:0] _t_pix_g;
reg  [7:0] _t_pix_b;

reg  [15:0] _d_cur_inv_y;
reg  [15:0] _q_cur_inv_y;
reg  [15:0] _d_pos_u;
reg  [15:0] _q_pos_u;
reg  [15:0] _d_pos_v;
reg  [15:0] _q_pos_v;
reg  [6:0] _d_lum;
reg  [6:0] _q_lum;
reg signed [15:0] _d__div_inum;
reg signed [15:0] _q__div_inum;
reg signed [15:0] _d__div_iden;
reg signed [15:0] _q__div_iden;
reg  [2:0] _d__idx_fsm0,_q__idx_fsm0;
reg  _autorun = 0;
reg  _div_run = 0;
assign out_pix_r = _t_pix_r;
assign out_pix_g = _t_pix_g;
assign out_pix_b = _t_pix_b;
assign out_done = (_q__idx_fsm0 == 0) && _autorun
;
M_div16_M_frame_display_div div (
.in_inum(_q__div_inum),
.in_iden(_q__div_iden),
.out_ret(_w_div_ret),
.out_done(_w_div_done),
.in_run(_div_run),
.reset(reset),
.clock(clock));



`ifdef FORMAL
initial begin
assume(reset);
end
assume property($initstate || (out_done));
`endif
always @* begin
_d_cur_inv_y = _q_cur_inv_y;
_d_pos_u = _q_pos_u;
_d_pos_v = _q_pos_v;
_d_lum = _q_lum;
_d__div_inum = _q__div_inum;
_d__div_iden = _q__div_iden;
_d__idx_fsm0 = _q__idx_fsm0;
_div_run = 1;
_t_offs_y = 0;
_t_u = 0;
_t_v = 0;
_t_floor = 0;
// _always_pre
_t_pix_r = 0;

_t_pix_g = 0;

_t_pix_b = 0;

(* full_case *)
case (_q__idx_fsm0)
1: begin
// _top
_d__idx_fsm0 = 2;
end
2: begin
// __while__block_1
if (1) begin
// __block_2
// __block_4
_d__idx_fsm0 = 3;
end else begin
// __block_3
_d__idx_fsm0 = 0;
end
end
3: begin
// __while__block_5
if (in_pix_vblank==0) begin
// __block_6
// __block_8
if (in_pix_active) begin
// __block_9
// __block_11
if (in_pix_y<240) begin
// __block_12
// __block_14
_t_offs_y = 272-in_pix_y;

_t_floor = 0;

// __block_15
end else begin
// __block_13
// __block_16
_t_offs_y = in_pix_y-208;

_t_floor = 1;

// __block_17
end
// 'after'
// __block_18
if (_t_offs_y>=35&&_t_offs_y<200) begin
// __block_19
// __block_21
if (in_pix_x==0) begin
// __block_22
// __block_24
_d_cur_inv_y = _w_div_ret;

if (_d_cur_inv_y[3+:7]<=70) begin
// __block_25
// __block_27
_d_lum = 70-_d_cur_inv_y[3+:7];

if (_d_lum>63) begin
// __block_28
// __block_30
_d_lum = 63;

// __block_31
end else begin
// __block_29
end
// 'after'
// __block_32
// __block_33
end else begin
// __block_26
// __block_34
_d_lum = 0;

// __block_35
end
// 'after'
// __block_36

_d__div_inum = _c_maxv;
_d__div_iden = _t_offs_y;
_div_run = 0;
// __block_37
end else begin
// __block_23
end
// 'after'
// __block_38
_t_u = _q_pos_u+((in_pix_x-320)*_d_cur_inv_y)>>8;

_t_v = _q_pos_v+_d_cur_inv_y[0+:6];

if (_t_u[5+:1]^_t_v[5+:1]) begin
// __block_39
// __block_41
if (_t_u[4+:1]^_t_v[4+:1]) begin
// __block_42
// __block_44
_t_pix_r = _d_lum<<2;

_t_pix_g = _d_lum<<2;

_t_pix_b = _d_lum<<2;

// __block_45
end else begin
// __block_43
// __block_46
_t_pix_r = _d_lum[1+:6]<<2;

_t_pix_g = _d_lum[1+:6]<<2;

_t_pix_b = _d_lum[1+:6]<<2;

// __block_47
end
// 'after'
// __block_48
// __block_49
end else begin
// __block_40
// __block_50
if (_t_u[4+:1]^_t_v[4+:1]) begin
// __block_51
// __block_53
if (_t_floor) begin
// __block_54
// __block_56
_t_pix_g = _d_lum<<2;

// __block_57
end else begin
// __block_55
// __block_58
_t_pix_b = _d_lum<<2;

// __block_59
end
// 'after'
// __block_60
// __block_61
end else begin
// __block_52
// __block_62
if (_t_floor) begin
// __block_63
// __block_65
_t_pix_g = _d_lum[1+:6]<<2;

// __block_66
end else begin
// __block_64
// __block_67
_t_pix_b = _d_lum[1+:6]<<2;

// __block_68
end
// 'after'
// __block_69
// __block_70
end
// 'after'
// __block_71
// __block_72
end
// 'after'
// __block_73
// __block_74
end else begin
// __block_20
end
// 'after'
// __block_75
// __block_76
end else begin
// __block_10
end
// 'after'
// __block_77
// __block_78
_d__idx_fsm0 = 3;
end else begin
// __block_7
_d_pos_u = _q_pos_u+1024;

_d_pos_v = _q_pos_v+3;

_d__idx_fsm0 = 4;
end
end
4: begin
// __while__block_79
if (in_pix_vblank==1) begin
// __block_80
// __block_82
// __block_83
_d__idx_fsm0 = 4;
end else begin
// __block_81
// __block_84
_d__idx_fsm0 = 2;
end
end
0: begin 
end
default: begin 
_d__idx_fsm0 = {3{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// _always_post
// pipeline stage triggers
end

always @(posedge clock) begin
_q_cur_inv_y <= (reset) ? 0 : _d_cur_inv_y;
_q_pos_u <= (reset) ? 0 : _d_pos_u;
_q_pos_v <= (reset) ? 0 : _d_pos_v;
_q_lum <= (reset) ? 0 : _d_lum;
_q__div_inum <= _d__div_inum;
_q__div_iden <= _d__div_iden;
_q__idx_fsm0 <= reset ? 0 : ( ~_autorun ? 1 : _d__idx_fsm0);
_autorun <= reset ? 0 : 1;
end

endmodule


/*
[Bare framework] Leave empty, this is used when exporting to verilog
*/

// SL 2019, MIT license
module M_frame_display__mem_cos(
input      [1-1:0]             in_wenable0,
input      signed [24-1:0]     in_wdata0,
input      [9-1:0]                in_addr0,
input      [1-1:0]             in_wenable1,
input      [24-1:0]                 in_wdata1,
input      [9-1:0]                in_addr1,
output reg signed [24-1:0]     out_rdata0,
output reg signed [24-1:0]     out_rdata1,
input      clock0,
input      clock1
);
(* no_rw_check *) reg signed [24-1:0] buffer[512-1:0];
always @(posedge clock0) begin
  if (in_wenable0) begin
    buffer[in_addr0] <= in_wdata0;
  end else begin
    out_rdata0 <= buffer[in_addr0];
  end
end
always @(posedge clock1) begin
  if (in_wenable1) begin
    buffer[in_addr1] <= in_wdata1;
  end else begin
    out_rdata1 <= buffer[in_addr1];
  end
end
initial begin
 buffer[0] = 1024;
 buffer[1] = 1023;
 buffer[2] = 1023;
 buffer[3] = 1023;
 buffer[4] = 1022;
 buffer[5] = 1022;
 buffer[6] = 1021;
 buffer[7] = 1020;
 buffer[8] = 1019;
 buffer[9] = 1017;
 buffer[10] = 1016;
 buffer[11] = 1014;
 buffer[12] = 1012;
 buffer[13] = 1010;
 buffer[14] = 1008;
 buffer[15] = 1006;
 buffer[16] = 1004;
 buffer[17] = 1001;
 buffer[18] = 999;
 buffer[19] = 996;
 buffer[20] = 993;
 buffer[21] = 990;
 buffer[22] = 986;
 buffer[23] = 983;
 buffer[24] = 979;
 buffer[25] = 976;
 buffer[26] = 972;
 buffer[27] = 968;
 buffer[28] = 964;
 buffer[29] = 959;
 buffer[30] = 955;
 buffer[31] = 950;
 buffer[32] = 946;
 buffer[33] = 941;
 buffer[34] = 936;
 buffer[35] = 930;
 buffer[36] = 925;
 buffer[37] = 920;
 buffer[38] = 914;
 buffer[39] = 908;
 buffer[40] = 903;
 buffer[41] = 897;
 buffer[42] = 890;
 buffer[43] = 884;
 buffer[44] = 878;
 buffer[45] = 871;
 buffer[46] = 865;
 buffer[47] = 858;
 buffer[48] = 851;
 buffer[49] = 844;
 buffer[50] = 837;
 buffer[51] = 829;
 buffer[52] = 822;
 buffer[53] = 814;
 buffer[54] = 807;
 buffer[55] = 799;
 buffer[56] = 791;
 buffer[57] = 783;
 buffer[58] = 775;
 buffer[59] = 767;
 buffer[60] = 758;
 buffer[61] = 750;
 buffer[62] = 741;
 buffer[63] = 732;
 buffer[64] = 724;
 buffer[65] = 715;
 buffer[66] = 706;
 buffer[67] = 696;
 buffer[68] = 687;
 buffer[69] = 678;
 buffer[70] = 668;
 buffer[71] = 659;
 buffer[72] = 649;
 buffer[73] = 639;
 buffer[74] = 629;
 buffer[75] = 620;
 buffer[76] = 609;
 buffer[77] = 599;
 buffer[78] = 589;
 buffer[79] = 579;
 buffer[80] = 568;
 buffer[81] = 558;
 buffer[82] = 547;
 buffer[83] = 537;
 buffer[84] = 526;
 buffer[85] = 515;
 buffer[86] = 504;
 buffer[87] = 493;
 buffer[88] = 482;
 buffer[89] = 471;
 buffer[90] = 460;
 buffer[91] = 449;
 buffer[92] = 437;
 buffer[93] = 426;
 buffer[94] = 414;
 buffer[95] = 403;
 buffer[96] = 391;
 buffer[97] = 380;
 buffer[98] = 368;
 buffer[99] = 356;
 buffer[100] = 344;
 buffer[101] = 333;
 buffer[102] = 321;
 buffer[103] = 309;
 buffer[104] = 297;
 buffer[105] = 285;
 buffer[106] = 273;
 buffer[107] = 260;
 buffer[108] = 248;
 buffer[109] = 236;
 buffer[110] = 224;
 buffer[111] = 212;
 buffer[112] = 199;
 buffer[113] = 187;
 buffer[114] = 175;
 buffer[115] = 162;
 buffer[116] = 150;
 buffer[117] = 137;
 buffer[118] = 125;
 buffer[119] = 112;
 buffer[120] = 100;
 buffer[121] = 87;
 buffer[122] = 75;
 buffer[123] = 62;
 buffer[124] = 50;
 buffer[125] = 37;
 buffer[126] = 25;
 buffer[127] = 12;
 buffer[128] = 0;
 buffer[129] = -13;
 buffer[130] = -26;
 buffer[131] = -38;
 buffer[132] = -51;
 buffer[133] = -63;
 buffer[134] = -76;
 buffer[135] = -88;
 buffer[136] = -101;
 buffer[137] = -113;
 buffer[138] = -126;
 buffer[139] = -138;
 buffer[140] = -151;
 buffer[141] = -163;
 buffer[142] = -176;
 buffer[143] = -188;
 buffer[144] = -200;
 buffer[145] = -213;
 buffer[146] = -225;
 buffer[147] = -237;
 buffer[148] = -249;
 buffer[149] = -261;
 buffer[150] = -274;
 buffer[151] = -286;
 buffer[152] = -298;
 buffer[153] = -310;
 buffer[154] = -322;
 buffer[155] = -334;
 buffer[156] = -345;
 buffer[157] = -357;
 buffer[158] = -369;
 buffer[159] = -381;
 buffer[160] = -392;
 buffer[161] = -404;
 buffer[162] = -415;
 buffer[163] = -427;
 buffer[164] = -438;
 buffer[165] = -450;
 buffer[166] = -461;
 buffer[167] = -472;
 buffer[168] = -483;
 buffer[169] = -494;
 buffer[170] = -505;
 buffer[171] = -516;
 buffer[172] = -527;
 buffer[173] = -538;
 buffer[174] = -548;
 buffer[175] = -559;
 buffer[176] = -569;
 buffer[177] = -580;
 buffer[178] = -590;
 buffer[179] = -600;
 buffer[180] = -610;
 buffer[181] = -621;
 buffer[182] = -630;
 buffer[183] = -640;
 buffer[184] = -650;
 buffer[185] = -660;
 buffer[186] = -669;
 buffer[187] = -679;
 buffer[188] = -688;
 buffer[189] = -697;
 buffer[190] = -707;
 buffer[191] = -716;
 buffer[192] = -725;
 buffer[193] = -733;
 buffer[194] = -742;
 buffer[195] = -751;
 buffer[196] = -759;
 buffer[197] = -768;
 buffer[198] = -776;
 buffer[199] = -784;
 buffer[200] = -792;
 buffer[201] = -800;
 buffer[202] = -808;
 buffer[203] = -815;
 buffer[204] = -823;
 buffer[205] = -830;
 buffer[206] = -838;
 buffer[207] = -845;
 buffer[208] = -852;
 buffer[209] = -859;
 buffer[210] = -866;
 buffer[211] = -872;
 buffer[212] = -879;
 buffer[213] = -885;
 buffer[214] = -891;
 buffer[215] = -898;
 buffer[216] = -904;
 buffer[217] = -909;
 buffer[218] = -915;
 buffer[219] = -921;
 buffer[220] = -926;
 buffer[221] = -931;
 buffer[222] = -937;
 buffer[223] = -942;
 buffer[224] = -947;
 buffer[225] = -951;
 buffer[226] = -956;
 buffer[227] = -960;
 buffer[228] = -965;
 buffer[229] = -969;
 buffer[230] = -973;
 buffer[231] = -977;
 buffer[232] = -980;
 buffer[233] = -984;
 buffer[234] = -987;
 buffer[235] = -991;
 buffer[236] = -994;
 buffer[237] = -997;
 buffer[238] = -1000;
 buffer[239] = -1002;
 buffer[240] = -1005;
 buffer[241] = -1007;
 buffer[242] = -1009;
 buffer[243] = -1011;
 buffer[244] = -1013;
 buffer[245] = -1015;
 buffer[246] = -1017;
 buffer[247] = -1018;
 buffer[248] = -1020;
 buffer[249] = -1021;
 buffer[250] = -1022;
 buffer[251] = -1023;
 buffer[252] = -1023;
 buffer[253] = -1024;
 buffer[254] = -1024;
 buffer[255] = -1024;
 buffer[256] = -1024;
 buffer[257] = -1024;
 buffer[258] = -1024;
 buffer[259] = -1024;
 buffer[260] = -1023;
 buffer[261] = -1023;
 buffer[262] = -1022;
 buffer[263] = -1021;
 buffer[264] = -1020;
 buffer[265] = -1018;
 buffer[266] = -1017;
 buffer[267] = -1015;
 buffer[268] = -1013;
 buffer[269] = -1011;
 buffer[270] = -1009;
 buffer[271] = -1007;
 buffer[272] = -1005;
 buffer[273] = -1002;
 buffer[274] = -1000;
 buffer[275] = -997;
 buffer[276] = -994;
 buffer[277] = -991;
 buffer[278] = -987;
 buffer[279] = -984;
 buffer[280] = -980;
 buffer[281] = -977;
 buffer[282] = -973;
 buffer[283] = -969;
 buffer[284] = -965;
 buffer[285] = -960;
 buffer[286] = -956;
 buffer[287] = -951;
 buffer[288] = -947;
 buffer[289] = -942;
 buffer[290] = -937;
 buffer[291] = -931;
 buffer[292] = -926;
 buffer[293] = -921;
 buffer[294] = -915;
 buffer[295] = -909;
 buffer[296] = -904;
 buffer[297] = -898;
 buffer[298] = -891;
 buffer[299] = -885;
 buffer[300] = -879;
 buffer[301] = -872;
 buffer[302] = -866;
 buffer[303] = -859;
 buffer[304] = -852;
 buffer[305] = -845;
 buffer[306] = -838;
 buffer[307] = -830;
 buffer[308] = -823;
 buffer[309] = -815;
 buffer[310] = -808;
 buffer[311] = -800;
 buffer[312] = -792;
 buffer[313] = -784;
 buffer[314] = -776;
 buffer[315] = -768;
 buffer[316] = -759;
 buffer[317] = -751;
 buffer[318] = -742;
 buffer[319] = -733;
 buffer[320] = -725;
 buffer[321] = -716;
 buffer[322] = -707;
 buffer[323] = -697;
 buffer[324] = -688;
 buffer[325] = -679;
 buffer[326] = -669;
 buffer[327] = -660;
 buffer[328] = -650;
 buffer[329] = -640;
 buffer[330] = -630;
 buffer[331] = -621;
 buffer[332] = -610;
 buffer[333] = -600;
 buffer[334] = -590;
 buffer[335] = -580;
 buffer[336] = -569;
 buffer[337] = -559;
 buffer[338] = -548;
 buffer[339] = -538;
 buffer[340] = -527;
 buffer[341] = -516;
 buffer[342] = -505;
 buffer[343] = -494;
 buffer[344] = -483;
 buffer[345] = -472;
 buffer[346] = -461;
 buffer[347] = -450;
 buffer[348] = -438;
 buffer[349] = -427;
 buffer[350] = -415;
 buffer[351] = -404;
 buffer[352] = -392;
 buffer[353] = -381;
 buffer[354] = -369;
 buffer[355] = -357;
 buffer[356] = -345;
 buffer[357] = -334;
 buffer[358] = -322;
 buffer[359] = -310;
 buffer[360] = -298;
 buffer[361] = -286;
 buffer[362] = -274;
 buffer[363] = -261;
 buffer[364] = -249;
 buffer[365] = -237;
 buffer[366] = -225;
 buffer[367] = -213;
 buffer[368] = -200;
 buffer[369] = -188;
 buffer[370] = -176;
 buffer[371] = -163;
 buffer[372] = -151;
 buffer[373] = -138;
 buffer[374] = -126;
 buffer[375] = -113;
 buffer[376] = -101;
 buffer[377] = -88;
 buffer[378] = -76;
 buffer[379] = -63;
 buffer[380] = -51;
 buffer[381] = -38;
 buffer[382] = -26;
 buffer[383] = -13;
 buffer[384] = -1;
 buffer[385] = 12;
 buffer[386] = 25;
 buffer[387] = 37;
 buffer[388] = 50;
 buffer[389] = 62;
 buffer[390] = 75;
 buffer[391] = 87;
 buffer[392] = 100;
 buffer[393] = 112;
 buffer[394] = 125;
 buffer[395] = 137;
 buffer[396] = 150;
 buffer[397] = 162;
 buffer[398] = 175;
 buffer[399] = 187;
 buffer[400] = 199;
 buffer[401] = 212;
 buffer[402] = 224;
 buffer[403] = 236;
 buffer[404] = 248;
 buffer[405] = 260;
 buffer[406] = 273;
 buffer[407] = 285;
 buffer[408] = 297;
 buffer[409] = 309;
 buffer[410] = 321;
 buffer[411] = 333;
 buffer[412] = 344;
 buffer[413] = 356;
 buffer[414] = 368;
 buffer[415] = 380;
 buffer[416] = 391;
 buffer[417] = 403;
 buffer[418] = 414;
 buffer[419] = 426;
 buffer[420] = 437;
 buffer[421] = 449;
 buffer[422] = 460;
 buffer[423] = 471;
 buffer[424] = 482;
 buffer[425] = 493;
 buffer[426] = 504;
 buffer[427] = 515;
 buffer[428] = 526;
 buffer[429] = 537;
 buffer[430] = 547;
 buffer[431] = 558;
 buffer[432] = 568;
 buffer[433] = 579;
 buffer[434] = 589;
 buffer[435] = 599;
 buffer[436] = 609;
 buffer[437] = 620;
 buffer[438] = 629;
 buffer[439] = 639;
 buffer[440] = 649;
 buffer[441] = 659;
 buffer[442] = 668;
 buffer[443] = 678;
 buffer[444] = 687;
 buffer[445] = 696;
 buffer[446] = 706;
 buffer[447] = 715;
 buffer[448] = 724;
 buffer[449] = 732;
 buffer[450] = 741;
 buffer[451] = 750;
 buffer[452] = 758;
 buffer[453] = 767;
 buffer[454] = 775;
 buffer[455] = 783;
 buffer[456] = 791;
 buffer[457] = 799;
 buffer[458] = 807;
 buffer[459] = 814;
 buffer[460] = 822;
 buffer[461] = 829;
 buffer[462] = 837;
 buffer[463] = 844;
 buffer[464] = 851;
 buffer[465] = 858;
 buffer[466] = 865;
 buffer[467] = 871;
 buffer[468] = 878;
 buffer[469] = 884;
 buffer[470] = 890;
 buffer[471] = 897;
 buffer[472] = 903;
 buffer[473] = 908;
 buffer[474] = 914;
 buffer[475] = 920;
 buffer[476] = 925;
 buffer[477] = 930;
 buffer[478] = 936;
 buffer[479] = 941;
 buffer[480] = 946;
 buffer[481] = 950;
 buffer[482] = 955;
 buffer[483] = 959;
 buffer[484] = 964;
 buffer[485] = 968;
 buffer[486] = 972;
 buffer[487] = 976;
 buffer[488] = 979;
 buffer[489] = 983;
 buffer[490] = 986;
 buffer[491] = 990;
 buffer[492] = 993;
 buffer[493] = 996;
 buffer[494] = 999;
 buffer[495] = 1001;
 buffer[496] = 1004;
 buffer[497] = 1006;
 buffer[498] = 1008;
 buffer[499] = 1010;
 buffer[500] = 1012;
 buffer[501] = 1014;
 buffer[502] = 1016;
 buffer[503] = 1017;
 buffer[504] = 1019;
 buffer[505] = 1020;
 buffer[506] = 1021;
 buffer[507] = 1022;
 buffer[508] = 1022;
 buffer[509] = 1023;
 buffer[510] = 1023;
 buffer[511] = 1023;
end

endmodule

// SL 2019, MIT license
module M_frame_display__mem_sin(
input      [1-1:0]             in_wenable0,
input      signed [24-1:0]     in_wdata0,
input      [9-1:0]                in_addr0,
input      [1-1:0]             in_wenable1,
input      [24-1:0]                 in_wdata1,
input      [9-1:0]                in_addr1,
output reg signed [24-1:0]     out_rdata0,
output reg signed [24-1:0]     out_rdata1,
input      clock0,
input      clock1
);
(* no_rw_check *) reg signed [24-1:0] buffer[512-1:0];
always @(posedge clock0) begin
  if (in_wenable0) begin
    buffer[in_addr0] <= in_wdata0;
  end else begin
    out_rdata0 <= buffer[in_addr0];
  end
end
always @(posedge clock1) begin
  if (in_wenable1) begin
    buffer[in_addr1] <= in_wdata1;
  end else begin
    out_rdata1 <= buffer[in_addr1];
  end
end
initial begin
 buffer[0] = 0;
 buffer[1] = 12;
 buffer[2] = 25;
 buffer[3] = 37;
 buffer[4] = 50;
 buffer[5] = 62;
 buffer[6] = 75;
 buffer[7] = 87;
 buffer[8] = 100;
 buffer[9] = 112;
 buffer[10] = 125;
 buffer[11] = 137;
 buffer[12] = 150;
 buffer[13] = 162;
 buffer[14] = 175;
 buffer[15] = 187;
 buffer[16] = 199;
 buffer[17] = 212;
 buffer[18] = 224;
 buffer[19] = 236;
 buffer[20] = 248;
 buffer[21] = 260;
 buffer[22] = 273;
 buffer[23] = 285;
 buffer[24] = 297;
 buffer[25] = 309;
 buffer[26] = 321;
 buffer[27] = 333;
 buffer[28] = 344;
 buffer[29] = 356;
 buffer[30] = 368;
 buffer[31] = 380;
 buffer[32] = 391;
 buffer[33] = 403;
 buffer[34] = 414;
 buffer[35] = 426;
 buffer[36] = 437;
 buffer[37] = 449;
 buffer[38] = 460;
 buffer[39] = 471;
 buffer[40] = 482;
 buffer[41] = 493;
 buffer[42] = 504;
 buffer[43] = 515;
 buffer[44] = 526;
 buffer[45] = 537;
 buffer[46] = 547;
 buffer[47] = 558;
 buffer[48] = 568;
 buffer[49] = 579;
 buffer[50] = 589;
 buffer[51] = 599;
 buffer[52] = 609;
 buffer[53] = 620;
 buffer[54] = 629;
 buffer[55] = 639;
 buffer[56] = 649;
 buffer[57] = 659;
 buffer[58] = 668;
 buffer[59] = 678;
 buffer[60] = 687;
 buffer[61] = 696;
 buffer[62] = 706;
 buffer[63] = 715;
 buffer[64] = 724;
 buffer[65] = 732;
 buffer[66] = 741;
 buffer[67] = 750;
 buffer[68] = 758;
 buffer[69] = 767;
 buffer[70] = 775;
 buffer[71] = 783;
 buffer[72] = 791;
 buffer[73] = 799;
 buffer[74] = 807;
 buffer[75] = 814;
 buffer[76] = 822;
 buffer[77] = 829;
 buffer[78] = 837;
 buffer[79] = 844;
 buffer[80] = 851;
 buffer[81] = 858;
 buffer[82] = 865;
 buffer[83] = 871;
 buffer[84] = 878;
 buffer[85] = 884;
 buffer[86] = 890;
 buffer[87] = 897;
 buffer[88] = 903;
 buffer[89] = 908;
 buffer[90] = 914;
 buffer[91] = 920;
 buffer[92] = 925;
 buffer[93] = 930;
 buffer[94] = 936;
 buffer[95] = 941;
 buffer[96] = 946;
 buffer[97] = 950;
 buffer[98] = 955;
 buffer[99] = 959;
 buffer[100] = 964;
 buffer[101] = 968;
 buffer[102] = 972;
 buffer[103] = 976;
 buffer[104] = 979;
 buffer[105] = 983;
 buffer[106] = 986;
 buffer[107] = 990;
 buffer[108] = 993;
 buffer[109] = 996;
 buffer[110] = 999;
 buffer[111] = 1001;
 buffer[112] = 1004;
 buffer[113] = 1006;
 buffer[114] = 1008;
 buffer[115] = 1010;
 buffer[116] = 1012;
 buffer[117] = 1014;
 buffer[118] = 1016;
 buffer[119] = 1017;
 buffer[120] = 1019;
 buffer[121] = 1020;
 buffer[122] = 1021;
 buffer[123] = 1022;
 buffer[124] = 1022;
 buffer[125] = 1023;
 buffer[126] = 1023;
 buffer[127] = 1023;
 buffer[128] = 1024;
 buffer[129] = 1023;
 buffer[130] = 1023;
 buffer[131] = 1023;
 buffer[132] = 1022;
 buffer[133] = 1022;
 buffer[134] = 1021;
 buffer[135] = 1020;
 buffer[136] = 1019;
 buffer[137] = 1017;
 buffer[138] = 1016;
 buffer[139] = 1014;
 buffer[140] = 1012;
 buffer[141] = 1010;
 buffer[142] = 1008;
 buffer[143] = 1006;
 buffer[144] = 1004;
 buffer[145] = 1001;
 buffer[146] = 999;
 buffer[147] = 996;
 buffer[148] = 993;
 buffer[149] = 990;
 buffer[150] = 986;
 buffer[151] = 983;
 buffer[152] = 979;
 buffer[153] = 976;
 buffer[154] = 972;
 buffer[155] = 968;
 buffer[156] = 964;
 buffer[157] = 959;
 buffer[158] = 955;
 buffer[159] = 950;
 buffer[160] = 946;
 buffer[161] = 941;
 buffer[162] = 936;
 buffer[163] = 930;
 buffer[164] = 925;
 buffer[165] = 920;
 buffer[166] = 914;
 buffer[167] = 908;
 buffer[168] = 903;
 buffer[169] = 897;
 buffer[170] = 890;
 buffer[171] = 884;
 buffer[172] = 878;
 buffer[173] = 871;
 buffer[174] = 865;
 buffer[175] = 858;
 buffer[176] = 851;
 buffer[177] = 844;
 buffer[178] = 837;
 buffer[179] = 829;
 buffer[180] = 822;
 buffer[181] = 814;
 buffer[182] = 807;
 buffer[183] = 799;
 buffer[184] = 791;
 buffer[185] = 783;
 buffer[186] = 775;
 buffer[187] = 767;
 buffer[188] = 758;
 buffer[189] = 750;
 buffer[190] = 741;
 buffer[191] = 732;
 buffer[192] = 724;
 buffer[193] = 715;
 buffer[194] = 706;
 buffer[195] = 696;
 buffer[196] = 687;
 buffer[197] = 678;
 buffer[198] = 668;
 buffer[199] = 659;
 buffer[200] = 649;
 buffer[201] = 639;
 buffer[202] = 629;
 buffer[203] = 620;
 buffer[204] = 609;
 buffer[205] = 599;
 buffer[206] = 589;
 buffer[207] = 579;
 buffer[208] = 568;
 buffer[209] = 558;
 buffer[210] = 547;
 buffer[211] = 537;
 buffer[212] = 526;
 buffer[213] = 515;
 buffer[214] = 504;
 buffer[215] = 493;
 buffer[216] = 482;
 buffer[217] = 471;
 buffer[218] = 460;
 buffer[219] = 449;
 buffer[220] = 437;
 buffer[221] = 426;
 buffer[222] = 414;
 buffer[223] = 403;
 buffer[224] = 391;
 buffer[225] = 380;
 buffer[226] = 368;
 buffer[227] = 356;
 buffer[228] = 344;
 buffer[229] = 333;
 buffer[230] = 321;
 buffer[231] = 309;
 buffer[232] = 297;
 buffer[233] = 285;
 buffer[234] = 273;
 buffer[235] = 260;
 buffer[236] = 248;
 buffer[237] = 236;
 buffer[238] = 224;
 buffer[239] = 212;
 buffer[240] = 199;
 buffer[241] = 187;
 buffer[242] = 175;
 buffer[243] = 162;
 buffer[244] = 150;
 buffer[245] = 137;
 buffer[246] = 125;
 buffer[247] = 112;
 buffer[248] = 100;
 buffer[249] = 87;
 buffer[250] = 75;
 buffer[251] = 62;
 buffer[252] = 50;
 buffer[253] = 37;
 buffer[254] = 25;
 buffer[255] = 12;
 buffer[256] = 0;
 buffer[257] = -13;
 buffer[258] = -26;
 buffer[259] = -38;
 buffer[260] = -51;
 buffer[261] = -63;
 buffer[262] = -76;
 buffer[263] = -88;
 buffer[264] = -101;
 buffer[265] = -113;
 buffer[266] = -126;
 buffer[267] = -138;
 buffer[268] = -151;
 buffer[269] = -163;
 buffer[270] = -176;
 buffer[271] = -188;
 buffer[272] = -200;
 buffer[273] = -213;
 buffer[274] = -225;
 buffer[275] = -237;
 buffer[276] = -249;
 buffer[277] = -261;
 buffer[278] = -274;
 buffer[279] = -286;
 buffer[280] = -298;
 buffer[281] = -310;
 buffer[282] = -322;
 buffer[283] = -334;
 buffer[284] = -345;
 buffer[285] = -357;
 buffer[286] = -369;
 buffer[287] = -381;
 buffer[288] = -392;
 buffer[289] = -404;
 buffer[290] = -415;
 buffer[291] = -427;
 buffer[292] = -438;
 buffer[293] = -450;
 buffer[294] = -461;
 buffer[295] = -472;
 buffer[296] = -483;
 buffer[297] = -494;
 buffer[298] = -505;
 buffer[299] = -516;
 buffer[300] = -527;
 buffer[301] = -538;
 buffer[302] = -548;
 buffer[303] = -559;
 buffer[304] = -569;
 buffer[305] = -580;
 buffer[306] = -590;
 buffer[307] = -600;
 buffer[308] = -610;
 buffer[309] = -621;
 buffer[310] = -630;
 buffer[311] = -640;
 buffer[312] = -650;
 buffer[313] = -660;
 buffer[314] = -669;
 buffer[315] = -679;
 buffer[316] = -688;
 buffer[317] = -697;
 buffer[318] = -707;
 buffer[319] = -716;
 buffer[320] = -725;
 buffer[321] = -733;
 buffer[322] = -742;
 buffer[323] = -751;
 buffer[324] = -759;
 buffer[325] = -768;
 buffer[326] = -776;
 buffer[327] = -784;
 buffer[328] = -792;
 buffer[329] = -800;
 buffer[330] = -808;
 buffer[331] = -815;
 buffer[332] = -823;
 buffer[333] = -830;
 buffer[334] = -838;
 buffer[335] = -845;
 buffer[336] = -852;
 buffer[337] = -859;
 buffer[338] = -866;
 buffer[339] = -872;
 buffer[340] = -879;
 buffer[341] = -885;
 buffer[342] = -891;
 buffer[343] = -898;
 buffer[344] = -904;
 buffer[345] = -909;
 buffer[346] = -915;
 buffer[347] = -921;
 buffer[348] = -926;
 buffer[349] = -931;
 buffer[350] = -937;
 buffer[351] = -942;
 buffer[352] = -947;
 buffer[353] = -951;
 buffer[354] = -956;
 buffer[355] = -960;
 buffer[356] = -965;
 buffer[357] = -969;
 buffer[358] = -973;
 buffer[359] = -977;
 buffer[360] = -980;
 buffer[361] = -984;
 buffer[362] = -987;
 buffer[363] = -991;
 buffer[364] = -994;
 buffer[365] = -997;
 buffer[366] = -1000;
 buffer[367] = -1002;
 buffer[368] = -1005;
 buffer[369] = -1007;
 buffer[370] = -1009;
 buffer[371] = -1011;
 buffer[372] = -1013;
 buffer[373] = -1015;
 buffer[374] = -1017;
 buffer[375] = -1018;
 buffer[376] = -1020;
 buffer[377] = -1021;
 buffer[378] = -1022;
 buffer[379] = -1023;
 buffer[380] = -1023;
 buffer[381] = -1024;
 buffer[382] = -1024;
 buffer[383] = -1024;
 buffer[384] = -1024;
 buffer[385] = -1024;
 buffer[386] = -1024;
 buffer[387] = -1024;
 buffer[388] = -1023;
 buffer[389] = -1023;
 buffer[390] = -1022;
 buffer[391] = -1021;
 buffer[392] = -1020;
 buffer[393] = -1018;
 buffer[394] = -1017;
 buffer[395] = -1015;
 buffer[396] = -1013;
 buffer[397] = -1011;
 buffer[398] = -1009;
 buffer[399] = -1007;
 buffer[400] = -1005;
 buffer[401] = -1002;
 buffer[402] = -1000;
 buffer[403] = -997;
 buffer[404] = -994;
 buffer[405] = -991;
 buffer[406] = -987;
 buffer[407] = -984;
 buffer[408] = -980;
 buffer[409] = -977;
 buffer[410] = -973;
 buffer[411] = -969;
 buffer[412] = -965;
 buffer[413] = -960;
 buffer[414] = -956;
 buffer[415] = -951;
 buffer[416] = -947;
 buffer[417] = -942;
 buffer[418] = -937;
 buffer[419] = -931;
 buffer[420] = -926;
 buffer[421] = -921;
 buffer[422] = -915;
 buffer[423] = -909;
 buffer[424] = -904;
 buffer[425] = -898;
 buffer[426] = -891;
 buffer[427] = -885;
 buffer[428] = -879;
 buffer[429] = -872;
 buffer[430] = -866;
 buffer[431] = -859;
 buffer[432] = -852;
 buffer[433] = -845;
 buffer[434] = -838;
 buffer[435] = -830;
 buffer[436] = -823;
 buffer[437] = -815;
 buffer[438] = -808;
 buffer[439] = -800;
 buffer[440] = -792;
 buffer[441] = -784;
 buffer[442] = -776;
 buffer[443] = -768;
 buffer[444] = -759;
 buffer[445] = -751;
 buffer[446] = -742;
 buffer[447] = -733;
 buffer[448] = -725;
 buffer[449] = -716;
 buffer[450] = -707;
 buffer[451] = -697;
 buffer[452] = -688;
 buffer[453] = -679;
 buffer[454] = -669;
 buffer[455] = -660;
 buffer[456] = -650;
 buffer[457] = -640;
 buffer[458] = -630;
 buffer[459] = -621;
 buffer[460] = -610;
 buffer[461] = -600;
 buffer[462] = -590;
 buffer[463] = -580;
 buffer[464] = -569;
 buffer[465] = -559;
 buffer[466] = -548;
 buffer[467] = -538;
 buffer[468] = -527;
 buffer[469] = -516;
 buffer[470] = -505;
 buffer[471] = -494;
 buffer[472] = -483;
 buffer[473] = -472;
 buffer[474] = -461;
 buffer[475] = -450;
 buffer[476] = -438;
 buffer[477] = -427;
 buffer[478] = -415;
 buffer[479] = -404;
 buffer[480] = -392;
 buffer[481] = -381;
 buffer[482] = -369;
 buffer[483] = -357;
 buffer[484] = -345;
 buffer[485] = -334;
 buffer[486] = -322;
 buffer[487] = -310;
 buffer[488] = -298;
 buffer[489] = -286;
 buffer[490] = -274;
 buffer[491] = -261;
 buffer[492] = -249;
 buffer[493] = -237;
 buffer[494] = -225;
 buffer[495] = -213;
 buffer[496] = -200;
 buffer[497] = -188;
 buffer[498] = -176;
 buffer[499] = -163;
 buffer[500] = -151;
 buffer[501] = -138;
 buffer[502] = -126;
 buffer[503] = -113;
 buffer[504] = -101;
 buffer[505] = -88;
 buffer[506] = -76;
 buffer[507] = -63;
 buffer[508] = -51;
 buffer[509] = -38;
 buffer[510] = -26;
 buffer[511] = -13;
end

endmodule

// SL 2019, MIT license
module M_frame_display__mem_invA(
input      [1-1:0]             in_wenable0,
input       [18-1:0]     in_wdata0,
input      [11-1:0]                in_addr0,
input      [1-1:0]             in_wenable1,
input      [18-1:0]                 in_wdata1,
input      [11-1:0]                in_addr1,
output reg  [18-1:0]     out_rdata0,
output reg  [18-1:0]     out_rdata1,
input      clock0,
input      clock1
);
(* no_rw_check *) reg  [18-1:0] buffer[2048-1:0];
always @(posedge clock0) begin
  if (in_wenable0) begin
    buffer[in_addr0] <= in_wdata0;
  end else begin
    out_rdata0 <= buffer[in_addr0];
  end
end
always @(posedge clock1) begin
  if (in_wenable1) begin
    buffer[in_addr1] <= in_wdata1;
  end else begin
    out_rdata1 <= buffer[in_addr1];
  end
end
initial begin
 buffer[0] = 131071;
 buffer[1] = 131071;
 buffer[2] = 131071;
 buffer[3] = 87381;
 buffer[4] = 65536;
 buffer[5] = 52428;
 buffer[6] = 43690;
 buffer[7] = 37449;
 buffer[8] = 32768;
 buffer[9] = 29127;
 buffer[10] = 26214;
 buffer[11] = 23831;
 buffer[12] = 21845;
 buffer[13] = 20164;
 buffer[14] = 18724;
 buffer[15] = 17476;
 buffer[16] = 16384;
 buffer[17] = 15420;
 buffer[18] = 14563;
 buffer[19] = 13797;
 buffer[20] = 13107;
 buffer[21] = 12483;
 buffer[22] = 11915;
 buffer[23] = 11397;
 buffer[24] = 10922;
 buffer[25] = 10485;
 buffer[26] = 10082;
 buffer[27] = 9709;
 buffer[28] = 9362;
 buffer[29] = 9039;
 buffer[30] = 8738;
 buffer[31] = 8456;
 buffer[32] = 8192;
 buffer[33] = 7943;
 buffer[34] = 7710;
 buffer[35] = 7489;
 buffer[36] = 7281;
 buffer[37] = 7084;
 buffer[38] = 6898;
 buffer[39] = 6721;
 buffer[40] = 6553;
 buffer[41] = 6393;
 buffer[42] = 6241;
 buffer[43] = 6096;
 buffer[44] = 5957;
 buffer[45] = 5825;
 buffer[46] = 5698;
 buffer[47] = 5577;
 buffer[48] = 5461;
 buffer[49] = 5349;
 buffer[50] = 5242;
 buffer[51] = 5140;
 buffer[52] = 5041;
 buffer[53] = 4946;
 buffer[54] = 4854;
 buffer[55] = 4766;
 buffer[56] = 4681;
 buffer[57] = 4599;
 buffer[58] = 4519;
 buffer[59] = 4443;
 buffer[60] = 4369;
 buffer[61] = 4297;
 buffer[62] = 4228;
 buffer[63] = 4161;
 buffer[64] = 4096;
 buffer[65] = 4032;
 buffer[66] = 3971;
 buffer[67] = 3912;
 buffer[68] = 3855;
 buffer[69] = 3799;
 buffer[70] = 3744;
 buffer[71] = 3692;
 buffer[72] = 3640;
 buffer[73] = 3591;
 buffer[74] = 3542;
 buffer[75] = 3495;
 buffer[76] = 3449;
 buffer[77] = 3404;
 buffer[78] = 3360;
 buffer[79] = 3318;
 buffer[80] = 3276;
 buffer[81] = 3236;
 buffer[82] = 3196;
 buffer[83] = 3158;
 buffer[84] = 3120;
 buffer[85] = 3084;
 buffer[86] = 3048;
 buffer[87] = 3013;
 buffer[88] = 2978;
 buffer[89] = 2945;
 buffer[90] = 2912;
 buffer[91] = 2880;
 buffer[92] = 2849;
 buffer[93] = 2818;
 buffer[94] = 2788;
 buffer[95] = 2759;
 buffer[96] = 2730;
 buffer[97] = 2702;
 buffer[98] = 2674;
 buffer[99] = 2647;
 buffer[100] = 2621;
 buffer[101] = 2595;
 buffer[102] = 2570;
 buffer[103] = 2545;
 buffer[104] = 2520;
 buffer[105] = 2496;
 buffer[106] = 2473;
 buffer[107] = 2449;
 buffer[108] = 2427;
 buffer[109] = 2404;
 buffer[110] = 2383;
 buffer[111] = 2361;
 buffer[112] = 2340;
 buffer[113] = 2319;
 buffer[114] = 2299;
 buffer[115] = 2279;
 buffer[116] = 2259;
 buffer[117] = 2240;
 buffer[118] = 2221;
 buffer[119] = 2202;
 buffer[120] = 2184;
 buffer[121] = 2166;
 buffer[122] = 2148;
 buffer[123] = 2131;
 buffer[124] = 2114;
 buffer[125] = 2097;
 buffer[126] = 2080;
 buffer[127] = 2064;
 buffer[128] = 2048;
 buffer[129] = 2032;
 buffer[130] = 2016;
 buffer[131] = 2001;
 buffer[132] = 1985;
 buffer[133] = 1971;
 buffer[134] = 1956;
 buffer[135] = 1941;
 buffer[136] = 1927;
 buffer[137] = 1913;
 buffer[138] = 1899;
 buffer[139] = 1885;
 buffer[140] = 1872;
 buffer[141] = 1859;
 buffer[142] = 1846;
 buffer[143] = 1833;
 buffer[144] = 1820;
 buffer[145] = 1807;
 buffer[146] = 1795;
 buffer[147] = 1783;
 buffer[148] = 1771;
 buffer[149] = 1759;
 buffer[150] = 1747;
 buffer[151] = 1736;
 buffer[152] = 1724;
 buffer[153] = 1713;
 buffer[154] = 1702;
 buffer[155] = 1691;
 buffer[156] = 1680;
 buffer[157] = 1669;
 buffer[158] = 1659;
 buffer[159] = 1648;
 buffer[160] = 1638;
 buffer[161] = 1628;
 buffer[162] = 1618;
 buffer[163] = 1608;
 buffer[164] = 1598;
 buffer[165] = 1588;
 buffer[166] = 1579;
 buffer[167] = 1569;
 buffer[168] = 1560;
 buffer[169] = 1551;
 buffer[170] = 1542;
 buffer[171] = 1533;
 buffer[172] = 1524;
 buffer[173] = 1515;
 buffer[174] = 1506;
 buffer[175] = 1497;
 buffer[176] = 1489;
 buffer[177] = 1481;
 buffer[178] = 1472;
 buffer[179] = 1464;
 buffer[180] = 1456;
 buffer[181] = 1448;
 buffer[182] = 1440;
 buffer[183] = 1432;
 buffer[184] = 1424;
 buffer[185] = 1416;
 buffer[186] = 1409;
 buffer[187] = 1401;
 buffer[188] = 1394;
 buffer[189] = 1387;
 buffer[190] = 1379;
 buffer[191] = 1372;
 buffer[192] = 1365;
 buffer[193] = 1358;
 buffer[194] = 1351;
 buffer[195] = 1344;
 buffer[196] = 1337;
 buffer[197] = 1330;
 buffer[198] = 1323;
 buffer[199] = 1317;
 buffer[200] = 1310;
 buffer[201] = 1304;
 buffer[202] = 1297;
 buffer[203] = 1291;
 buffer[204] = 1285;
 buffer[205] = 1278;
 buffer[206] = 1272;
 buffer[207] = 1266;
 buffer[208] = 1260;
 buffer[209] = 1254;
 buffer[210] = 1248;
 buffer[211] = 1242;
 buffer[212] = 1236;
 buffer[213] = 1230;
 buffer[214] = 1224;
 buffer[215] = 1219;
 buffer[216] = 1213;
 buffer[217] = 1208;
 buffer[218] = 1202;
 buffer[219] = 1197;
 buffer[220] = 1191;
 buffer[221] = 1186;
 buffer[222] = 1180;
 buffer[223] = 1175;
 buffer[224] = 1170;
 buffer[225] = 1165;
 buffer[226] = 1159;
 buffer[227] = 1154;
 buffer[228] = 1149;
 buffer[229] = 1144;
 buffer[230] = 1139;
 buffer[231] = 1134;
 buffer[232] = 1129;
 buffer[233] = 1125;
 buffer[234] = 1120;
 buffer[235] = 1115;
 buffer[236] = 1110;
 buffer[237] = 1106;
 buffer[238] = 1101;
 buffer[239] = 1096;
 buffer[240] = 1092;
 buffer[241] = 1087;
 buffer[242] = 1083;
 buffer[243] = 1078;
 buffer[244] = 1074;
 buffer[245] = 1069;
 buffer[246] = 1065;
 buffer[247] = 1061;
 buffer[248] = 1057;
 buffer[249] = 1052;
 buffer[250] = 1048;
 buffer[251] = 1044;
 buffer[252] = 1040;
 buffer[253] = 1036;
 buffer[254] = 1032;
 buffer[255] = 1028;
 buffer[256] = 1024;
 buffer[257] = 1020;
 buffer[258] = 1016;
 buffer[259] = 1012;
 buffer[260] = 1008;
 buffer[261] = 1004;
 buffer[262] = 1000;
 buffer[263] = 996;
 buffer[264] = 992;
 buffer[265] = 989;
 buffer[266] = 985;
 buffer[267] = 981;
 buffer[268] = 978;
 buffer[269] = 974;
 buffer[270] = 970;
 buffer[271] = 967;
 buffer[272] = 963;
 buffer[273] = 960;
 buffer[274] = 956;
 buffer[275] = 953;
 buffer[276] = 949;
 buffer[277] = 946;
 buffer[278] = 942;
 buffer[279] = 939;
 buffer[280] = 936;
 buffer[281] = 932;
 buffer[282] = 929;
 buffer[283] = 926;
 buffer[284] = 923;
 buffer[285] = 919;
 buffer[286] = 916;
 buffer[287] = 913;
 buffer[288] = 910;
 buffer[289] = 907;
 buffer[290] = 903;
 buffer[291] = 900;
 buffer[292] = 897;
 buffer[293] = 894;
 buffer[294] = 891;
 buffer[295] = 888;
 buffer[296] = 885;
 buffer[297] = 882;
 buffer[298] = 879;
 buffer[299] = 876;
 buffer[300] = 873;
 buffer[301] = 870;
 buffer[302] = 868;
 buffer[303] = 865;
 buffer[304] = 862;
 buffer[305] = 859;
 buffer[306] = 856;
 buffer[307] = 853;
 buffer[308] = 851;
 buffer[309] = 848;
 buffer[310] = 845;
 buffer[311] = 842;
 buffer[312] = 840;
 buffer[313] = 837;
 buffer[314] = 834;
 buffer[315] = 832;
 buffer[316] = 829;
 buffer[317] = 826;
 buffer[318] = 824;
 buffer[319] = 821;
 buffer[320] = 819;
 buffer[321] = 816;
 buffer[322] = 814;
 buffer[323] = 811;
 buffer[324] = 809;
 buffer[325] = 806;
 buffer[326] = 804;
 buffer[327] = 801;
 buffer[328] = 799;
 buffer[329] = 796;
 buffer[330] = 794;
 buffer[331] = 791;
 buffer[332] = 789;
 buffer[333] = 787;
 buffer[334] = 784;
 buffer[335] = 782;
 buffer[336] = 780;
 buffer[337] = 777;
 buffer[338] = 775;
 buffer[339] = 773;
 buffer[340] = 771;
 buffer[341] = 768;
 buffer[342] = 766;
 buffer[343] = 764;
 buffer[344] = 762;
 buffer[345] = 759;
 buffer[346] = 757;
 buffer[347] = 755;
 buffer[348] = 753;
 buffer[349] = 751;
 buffer[350] = 748;
 buffer[351] = 746;
 buffer[352] = 744;
 buffer[353] = 742;
 buffer[354] = 740;
 buffer[355] = 738;
 buffer[356] = 736;
 buffer[357] = 734;
 buffer[358] = 732;
 buffer[359] = 730;
 buffer[360] = 728;
 buffer[361] = 726;
 buffer[362] = 724;
 buffer[363] = 722;
 buffer[364] = 720;
 buffer[365] = 718;
 buffer[366] = 716;
 buffer[367] = 714;
 buffer[368] = 712;
 buffer[369] = 710;
 buffer[370] = 708;
 buffer[371] = 706;
 buffer[372] = 704;
 buffer[373] = 702;
 buffer[374] = 700;
 buffer[375] = 699;
 buffer[376] = 697;
 buffer[377] = 695;
 buffer[378] = 693;
 buffer[379] = 691;
 buffer[380] = 689;
 buffer[381] = 688;
 buffer[382] = 686;
 buffer[383] = 684;
 buffer[384] = 682;
 buffer[385] = 680;
 buffer[386] = 679;
 buffer[387] = 677;
 buffer[388] = 675;
 buffer[389] = 673;
 buffer[390] = 672;
 buffer[391] = 670;
 buffer[392] = 668;
 buffer[393] = 667;
 buffer[394] = 665;
 buffer[395] = 663;
 buffer[396] = 661;
 buffer[397] = 660;
 buffer[398] = 658;
 buffer[399] = 657;
 buffer[400] = 655;
 buffer[401] = 653;
 buffer[402] = 652;
 buffer[403] = 650;
 buffer[404] = 648;
 buffer[405] = 647;
 buffer[406] = 645;
 buffer[407] = 644;
 buffer[408] = 642;
 buffer[409] = 640;
 buffer[410] = 639;
 buffer[411] = 637;
 buffer[412] = 636;
 buffer[413] = 634;
 buffer[414] = 633;
 buffer[415] = 631;
 buffer[416] = 630;
 buffer[417] = 628;
 buffer[418] = 627;
 buffer[419] = 625;
 buffer[420] = 624;
 buffer[421] = 622;
 buffer[422] = 621;
 buffer[423] = 619;
 buffer[424] = 618;
 buffer[425] = 616;
 buffer[426] = 615;
 buffer[427] = 613;
 buffer[428] = 612;
 buffer[429] = 611;
 buffer[430] = 609;
 buffer[431] = 608;
 buffer[432] = 606;
 buffer[433] = 605;
 buffer[434] = 604;
 buffer[435] = 602;
 buffer[436] = 601;
 buffer[437] = 599;
 buffer[438] = 598;
 buffer[439] = 597;
 buffer[440] = 595;
 buffer[441] = 594;
 buffer[442] = 593;
 buffer[443] = 591;
 buffer[444] = 590;
 buffer[445] = 589;
 buffer[446] = 587;
 buffer[447] = 586;
 buffer[448] = 585;
 buffer[449] = 583;
 buffer[450] = 582;
 buffer[451] = 581;
 buffer[452] = 579;
 buffer[453] = 578;
 buffer[454] = 577;
 buffer[455] = 576;
 buffer[456] = 574;
 buffer[457] = 573;
 buffer[458] = 572;
 buffer[459] = 571;
 buffer[460] = 569;
 buffer[461] = 568;
 buffer[462] = 567;
 buffer[463] = 566;
 buffer[464] = 564;
 buffer[465] = 563;
 buffer[466] = 562;
 buffer[467] = 561;
 buffer[468] = 560;
 buffer[469] = 558;
 buffer[470] = 557;
 buffer[471] = 556;
 buffer[472] = 555;
 buffer[473] = 554;
 buffer[474] = 553;
 buffer[475] = 551;
 buffer[476] = 550;
 buffer[477] = 549;
 buffer[478] = 548;
 buffer[479] = 547;
 buffer[480] = 546;
 buffer[481] = 544;
 buffer[482] = 543;
 buffer[483] = 542;
 buffer[484] = 541;
 buffer[485] = 540;
 buffer[486] = 539;
 buffer[487] = 538;
 buffer[488] = 537;
 buffer[489] = 536;
 buffer[490] = 534;
 buffer[491] = 533;
 buffer[492] = 532;
 buffer[493] = 531;
 buffer[494] = 530;
 buffer[495] = 529;
 buffer[496] = 528;
 buffer[497] = 527;
 buffer[498] = 526;
 buffer[499] = 525;
 buffer[500] = 524;
 buffer[501] = 523;
 buffer[502] = 522;
 buffer[503] = 521;
 buffer[504] = 520;
 buffer[505] = 519;
 buffer[506] = 518;
 buffer[507] = 517;
 buffer[508] = 516;
 buffer[509] = 515;
 buffer[510] = 514;
 buffer[511] = 513;
 buffer[512] = 512;
 buffer[513] = 511;
 buffer[514] = 510;
 buffer[515] = 509;
 buffer[516] = 508;
 buffer[517] = 507;
 buffer[518] = 506;
 buffer[519] = 505;
 buffer[520] = 504;
 buffer[521] = 503;
 buffer[522] = 502;
 buffer[523] = 501;
 buffer[524] = 500;
 buffer[525] = 499;
 buffer[526] = 498;
 buffer[527] = 497;
 buffer[528] = 496;
 buffer[529] = 495;
 buffer[530] = 494;
 buffer[531] = 493;
 buffer[532] = 492;
 buffer[533] = 491;
 buffer[534] = 490;
 buffer[535] = 489;
 buffer[536] = 489;
 buffer[537] = 488;
 buffer[538] = 487;
 buffer[539] = 486;
 buffer[540] = 485;
 buffer[541] = 484;
 buffer[542] = 483;
 buffer[543] = 482;
 buffer[544] = 481;
 buffer[545] = 480;
 buffer[546] = 480;
 buffer[547] = 479;
 buffer[548] = 478;
 buffer[549] = 477;
 buffer[550] = 476;
 buffer[551] = 475;
 buffer[552] = 474;
 buffer[553] = 474;
 buffer[554] = 473;
 buffer[555] = 472;
 buffer[556] = 471;
 buffer[557] = 470;
 buffer[558] = 469;
 buffer[559] = 468;
 buffer[560] = 468;
 buffer[561] = 467;
 buffer[562] = 466;
 buffer[563] = 465;
 buffer[564] = 464;
 buffer[565] = 463;
 buffer[566] = 463;
 buffer[567] = 462;
 buffer[568] = 461;
 buffer[569] = 460;
 buffer[570] = 459;
 buffer[571] = 459;
 buffer[572] = 458;
 buffer[573] = 457;
 buffer[574] = 456;
 buffer[575] = 455;
 buffer[576] = 455;
 buffer[577] = 454;
 buffer[578] = 453;
 buffer[579] = 452;
 buffer[580] = 451;
 buffer[581] = 451;
 buffer[582] = 450;
 buffer[583] = 449;
 buffer[584] = 448;
 buffer[585] = 448;
 buffer[586] = 447;
 buffer[587] = 446;
 buffer[588] = 445;
 buffer[589] = 445;
 buffer[590] = 444;
 buffer[591] = 443;
 buffer[592] = 442;
 buffer[593] = 442;
 buffer[594] = 441;
 buffer[595] = 440;
 buffer[596] = 439;
 buffer[597] = 439;
 buffer[598] = 438;
 buffer[599] = 437;
 buffer[600] = 436;
 buffer[601] = 436;
 buffer[602] = 435;
 buffer[603] = 434;
 buffer[604] = 434;
 buffer[605] = 433;
 buffer[606] = 432;
 buffer[607] = 431;
 buffer[608] = 431;
 buffer[609] = 430;
 buffer[610] = 429;
 buffer[611] = 429;
 buffer[612] = 428;
 buffer[613] = 427;
 buffer[614] = 426;
 buffer[615] = 426;
 buffer[616] = 425;
 buffer[617] = 424;
 buffer[618] = 424;
 buffer[619] = 423;
 buffer[620] = 422;
 buffer[621] = 422;
 buffer[622] = 421;
 buffer[623] = 420;
 buffer[624] = 420;
 buffer[625] = 419;
 buffer[626] = 418;
 buffer[627] = 418;
 buffer[628] = 417;
 buffer[629] = 416;
 buffer[630] = 416;
 buffer[631] = 415;
 buffer[632] = 414;
 buffer[633] = 414;
 buffer[634] = 413;
 buffer[635] = 412;
 buffer[636] = 412;
 buffer[637] = 411;
 buffer[638] = 410;
 buffer[639] = 410;
 buffer[640] = 409;
 buffer[641] = 408;
 buffer[642] = 408;
 buffer[643] = 407;
 buffer[644] = 407;
 buffer[645] = 406;
 buffer[646] = 405;
 buffer[647] = 405;
 buffer[648] = 404;
 buffer[649] = 403;
 buffer[650] = 403;
 buffer[651] = 402;
 buffer[652] = 402;
 buffer[653] = 401;
 buffer[654] = 400;
 buffer[655] = 400;
 buffer[656] = 399;
 buffer[657] = 399;
 buffer[658] = 398;
 buffer[659] = 397;
 buffer[660] = 397;
 buffer[661] = 396;
 buffer[662] = 395;
 buffer[663] = 395;
 buffer[664] = 394;
 buffer[665] = 394;
 buffer[666] = 393;
 buffer[667] = 393;
 buffer[668] = 392;
 buffer[669] = 391;
 buffer[670] = 391;
 buffer[671] = 390;
 buffer[672] = 390;
 buffer[673] = 389;
 buffer[674] = 388;
 buffer[675] = 388;
 buffer[676] = 387;
 buffer[677] = 387;
 buffer[678] = 386;
 buffer[679] = 386;
 buffer[680] = 385;
 buffer[681] = 384;
 buffer[682] = 384;
 buffer[683] = 383;
 buffer[684] = 383;
 buffer[685] = 382;
 buffer[686] = 382;
 buffer[687] = 381;
 buffer[688] = 381;
 buffer[689] = 380;
 buffer[690] = 379;
 buffer[691] = 379;
 buffer[692] = 378;
 buffer[693] = 378;
 buffer[694] = 377;
 buffer[695] = 377;
 buffer[696] = 376;
 buffer[697] = 376;
 buffer[698] = 375;
 buffer[699] = 375;
 buffer[700] = 374;
 buffer[701] = 373;
 buffer[702] = 373;
 buffer[703] = 372;
 buffer[704] = 372;
 buffer[705] = 371;
 buffer[706] = 371;
 buffer[707] = 370;
 buffer[708] = 370;
 buffer[709] = 369;
 buffer[710] = 369;
 buffer[711] = 368;
 buffer[712] = 368;
 buffer[713] = 367;
 buffer[714] = 367;
 buffer[715] = 366;
 buffer[716] = 366;
 buffer[717] = 365;
 buffer[718] = 365;
 buffer[719] = 364;
 buffer[720] = 364;
 buffer[721] = 363;
 buffer[722] = 363;
 buffer[723] = 362;
 buffer[724] = 362;
 buffer[725] = 361;
 buffer[726] = 361;
 buffer[727] = 360;
 buffer[728] = 360;
 buffer[729] = 359;
 buffer[730] = 359;
 buffer[731] = 358;
 buffer[732] = 358;
 buffer[733] = 357;
 buffer[734] = 357;
 buffer[735] = 356;
 buffer[736] = 356;
 buffer[737] = 355;
 buffer[738] = 355;
 buffer[739] = 354;
 buffer[740] = 354;
 buffer[741] = 353;
 buffer[742] = 353;
 buffer[743] = 352;
 buffer[744] = 352;
 buffer[745] = 351;
 buffer[746] = 351;
 buffer[747] = 350;
 buffer[748] = 350;
 buffer[749] = 349;
 buffer[750] = 349;
 buffer[751] = 349;
 buffer[752] = 348;
 buffer[753] = 348;
 buffer[754] = 347;
 buffer[755] = 347;
 buffer[756] = 346;
 buffer[757] = 346;
 buffer[758] = 345;
 buffer[759] = 345;
 buffer[760] = 344;
 buffer[761] = 344;
 buffer[762] = 344;
 buffer[763] = 343;
 buffer[764] = 343;
 buffer[765] = 342;
 buffer[766] = 342;
 buffer[767] = 341;
 buffer[768] = 341;
 buffer[769] = 340;
 buffer[770] = 340;
 buffer[771] = 340;
 buffer[772] = 339;
 buffer[773] = 339;
 buffer[774] = 338;
 buffer[775] = 338;
 buffer[776] = 337;
 buffer[777] = 337;
 buffer[778] = 336;
 buffer[779] = 336;
 buffer[780] = 336;
 buffer[781] = 335;
 buffer[782] = 335;
 buffer[783] = 334;
 buffer[784] = 334;
 buffer[785] = 333;
 buffer[786] = 333;
 buffer[787] = 333;
 buffer[788] = 332;
 buffer[789] = 332;
 buffer[790] = 331;
 buffer[791] = 331;
 buffer[792] = 330;
 buffer[793] = 330;
 buffer[794] = 330;
 buffer[795] = 329;
 buffer[796] = 329;
 buffer[797] = 328;
 buffer[798] = 328;
 buffer[799] = 328;
 buffer[800] = 327;
 buffer[801] = 327;
 buffer[802] = 326;
 buffer[803] = 326;
 buffer[804] = 326;
 buffer[805] = 325;
 buffer[806] = 325;
 buffer[807] = 324;
 buffer[808] = 324;
 buffer[809] = 324;
 buffer[810] = 323;
 buffer[811] = 323;
 buffer[812] = 322;
 buffer[813] = 322;
 buffer[814] = 322;
 buffer[815] = 321;
 buffer[816] = 321;
 buffer[817] = 320;
 buffer[818] = 320;
 buffer[819] = 320;
 buffer[820] = 319;
 buffer[821] = 319;
 buffer[822] = 318;
 buffer[823] = 318;
 buffer[824] = 318;
 buffer[825] = 317;
 buffer[826] = 317;
 buffer[827] = 316;
 buffer[828] = 316;
 buffer[829] = 316;
 buffer[830] = 315;
 buffer[831] = 315;
 buffer[832] = 315;
 buffer[833] = 314;
 buffer[834] = 314;
 buffer[835] = 313;
 buffer[836] = 313;
 buffer[837] = 313;
 buffer[838] = 312;
 buffer[839] = 312;
 buffer[840] = 312;
 buffer[841] = 311;
 buffer[842] = 311;
 buffer[843] = 310;
 buffer[844] = 310;
 buffer[845] = 310;
 buffer[846] = 309;
 buffer[847] = 309;
 buffer[848] = 309;
 buffer[849] = 308;
 buffer[850] = 308;
 buffer[851] = 308;
 buffer[852] = 307;
 buffer[853] = 307;
 buffer[854] = 306;
 buffer[855] = 306;
 buffer[856] = 306;
 buffer[857] = 305;
 buffer[858] = 305;
 buffer[859] = 305;
 buffer[860] = 304;
 buffer[861] = 304;
 buffer[862] = 304;
 buffer[863] = 303;
 buffer[864] = 303;
 buffer[865] = 303;
 buffer[866] = 302;
 buffer[867] = 302;
 buffer[868] = 302;
 buffer[869] = 301;
 buffer[870] = 301;
 buffer[871] = 300;
 buffer[872] = 300;
 buffer[873] = 300;
 buffer[874] = 299;
 buffer[875] = 299;
 buffer[876] = 299;
 buffer[877] = 298;
 buffer[878] = 298;
 buffer[879] = 298;
 buffer[880] = 297;
 buffer[881] = 297;
 buffer[882] = 297;
 buffer[883] = 296;
 buffer[884] = 296;
 buffer[885] = 296;
 buffer[886] = 295;
 buffer[887] = 295;
 buffer[888] = 295;
 buffer[889] = 294;
 buffer[890] = 294;
 buffer[891] = 294;
 buffer[892] = 293;
 buffer[893] = 293;
 buffer[894] = 293;
 buffer[895] = 292;
 buffer[896] = 292;
 buffer[897] = 292;
 buffer[898] = 291;
 buffer[899] = 291;
 buffer[900] = 291;
 buffer[901] = 290;
 buffer[902] = 290;
 buffer[903] = 290;
 buffer[904] = 289;
 buffer[905] = 289;
 buffer[906] = 289;
 buffer[907] = 289;
 buffer[908] = 288;
 buffer[909] = 288;
 buffer[910] = 288;
 buffer[911] = 287;
 buffer[912] = 287;
 buffer[913] = 287;
 buffer[914] = 286;
 buffer[915] = 286;
 buffer[916] = 286;
 buffer[917] = 285;
 buffer[918] = 285;
 buffer[919] = 285;
 buffer[920] = 284;
 buffer[921] = 284;
 buffer[922] = 284;
 buffer[923] = 284;
 buffer[924] = 283;
 buffer[925] = 283;
 buffer[926] = 283;
 buffer[927] = 282;
 buffer[928] = 282;
 buffer[929] = 282;
 buffer[930] = 281;
 buffer[931] = 281;
 buffer[932] = 281;
 buffer[933] = 280;
 buffer[934] = 280;
 buffer[935] = 280;
 buffer[936] = 280;
 buffer[937] = 279;
 buffer[938] = 279;
 buffer[939] = 279;
 buffer[940] = 278;
 buffer[941] = 278;
 buffer[942] = 278;
 buffer[943] = 277;
 buffer[944] = 277;
 buffer[945] = 277;
 buffer[946] = 277;
 buffer[947] = 276;
 buffer[948] = 276;
 buffer[949] = 276;
 buffer[950] = 275;
 buffer[951] = 275;
 buffer[952] = 275;
 buffer[953] = 275;
 buffer[954] = 274;
 buffer[955] = 274;
 buffer[956] = 274;
 buffer[957] = 273;
 buffer[958] = 273;
 buffer[959] = 273;
 buffer[960] = 273;
 buffer[961] = 272;
 buffer[962] = 272;
 buffer[963] = 272;
 buffer[964] = 271;
 buffer[965] = 271;
 buffer[966] = 271;
 buffer[967] = 271;
 buffer[968] = 270;
 buffer[969] = 270;
 buffer[970] = 270;
 buffer[971] = 269;
 buffer[972] = 269;
 buffer[973] = 269;
 buffer[974] = 269;
 buffer[975] = 268;
 buffer[976] = 268;
 buffer[977] = 268;
 buffer[978] = 268;
 buffer[979] = 267;
 buffer[980] = 267;
 buffer[981] = 267;
 buffer[982] = 266;
 buffer[983] = 266;
 buffer[984] = 266;
 buffer[985] = 266;
 buffer[986] = 265;
 buffer[987] = 265;
 buffer[988] = 265;
 buffer[989] = 265;
 buffer[990] = 264;
 buffer[991] = 264;
 buffer[992] = 264;
 buffer[993] = 263;
 buffer[994] = 263;
 buffer[995] = 263;
 buffer[996] = 263;
 buffer[997] = 262;
 buffer[998] = 262;
 buffer[999] = 262;
 buffer[1000] = 262;
 buffer[1001] = 261;
 buffer[1002] = 261;
 buffer[1003] = 261;
 buffer[1004] = 261;
 buffer[1005] = 260;
 buffer[1006] = 260;
 buffer[1007] = 260;
 buffer[1008] = 260;
 buffer[1009] = 259;
 buffer[1010] = 259;
 buffer[1011] = 259;
 buffer[1012] = 259;
 buffer[1013] = 258;
 buffer[1014] = 258;
 buffer[1015] = 258;
 buffer[1016] = 258;
 buffer[1017] = 257;
 buffer[1018] = 257;
 buffer[1019] = 257;
 buffer[1020] = 257;
 buffer[1021] = 256;
 buffer[1022] = 256;
 buffer[1023] = 256;
 buffer[1024] = 256;
 buffer[1025] = 255;
 buffer[1026] = 255;
 buffer[1027] = 255;
 buffer[1028] = 255;
 buffer[1029] = 254;
 buffer[1030] = 254;
 buffer[1031] = 254;
 buffer[1032] = 254;
 buffer[1033] = 253;
 buffer[1034] = 253;
 buffer[1035] = 253;
 buffer[1036] = 253;
 buffer[1037] = 252;
 buffer[1038] = 252;
 buffer[1039] = 252;
 buffer[1040] = 252;
 buffer[1041] = 251;
 buffer[1042] = 251;
 buffer[1043] = 251;
 buffer[1044] = 251;
 buffer[1045] = 250;
 buffer[1046] = 250;
 buffer[1047] = 250;
 buffer[1048] = 250;
 buffer[1049] = 249;
 buffer[1050] = 249;
 buffer[1051] = 249;
 buffer[1052] = 249;
 buffer[1053] = 248;
 buffer[1054] = 248;
 buffer[1055] = 248;
 buffer[1056] = 248;
 buffer[1057] = 248;
 buffer[1058] = 247;
 buffer[1059] = 247;
 buffer[1060] = 247;
 buffer[1061] = 247;
 buffer[1062] = 246;
 buffer[1063] = 246;
 buffer[1064] = 246;
 buffer[1065] = 246;
 buffer[1066] = 245;
 buffer[1067] = 245;
 buffer[1068] = 245;
 buffer[1069] = 245;
 buffer[1070] = 244;
 buffer[1071] = 244;
 buffer[1072] = 244;
 buffer[1073] = 244;
 buffer[1074] = 244;
 buffer[1075] = 243;
 buffer[1076] = 243;
 buffer[1077] = 243;
 buffer[1078] = 243;
 buffer[1079] = 242;
 buffer[1080] = 242;
 buffer[1081] = 242;
 buffer[1082] = 242;
 buffer[1083] = 242;
 buffer[1084] = 241;
 buffer[1085] = 241;
 buffer[1086] = 241;
 buffer[1087] = 241;
 buffer[1088] = 240;
 buffer[1089] = 240;
 buffer[1090] = 240;
 buffer[1091] = 240;
 buffer[1092] = 240;
 buffer[1093] = 239;
 buffer[1094] = 239;
 buffer[1095] = 239;
 buffer[1096] = 239;
 buffer[1097] = 238;
 buffer[1098] = 238;
 buffer[1099] = 238;
 buffer[1100] = 238;
 buffer[1101] = 238;
 buffer[1102] = 237;
 buffer[1103] = 237;
 buffer[1104] = 237;
 buffer[1105] = 237;
 buffer[1106] = 237;
 buffer[1107] = 236;
 buffer[1108] = 236;
 buffer[1109] = 236;
 buffer[1110] = 236;
 buffer[1111] = 235;
 buffer[1112] = 235;
 buffer[1113] = 235;
 buffer[1114] = 235;
 buffer[1115] = 235;
 buffer[1116] = 234;
 buffer[1117] = 234;
 buffer[1118] = 234;
 buffer[1119] = 234;
 buffer[1120] = 234;
 buffer[1121] = 233;
 buffer[1122] = 233;
 buffer[1123] = 233;
 buffer[1124] = 233;
 buffer[1125] = 233;
 buffer[1126] = 232;
 buffer[1127] = 232;
 buffer[1128] = 232;
 buffer[1129] = 232;
 buffer[1130] = 231;
 buffer[1131] = 231;
 buffer[1132] = 231;
 buffer[1133] = 231;
 buffer[1134] = 231;
 buffer[1135] = 230;
 buffer[1136] = 230;
 buffer[1137] = 230;
 buffer[1138] = 230;
 buffer[1139] = 230;
 buffer[1140] = 229;
 buffer[1141] = 229;
 buffer[1142] = 229;
 buffer[1143] = 229;
 buffer[1144] = 229;
 buffer[1145] = 228;
 buffer[1146] = 228;
 buffer[1147] = 228;
 buffer[1148] = 228;
 buffer[1149] = 228;
 buffer[1150] = 227;
 buffer[1151] = 227;
 buffer[1152] = 227;
 buffer[1153] = 227;
 buffer[1154] = 227;
 buffer[1155] = 226;
 buffer[1156] = 226;
 buffer[1157] = 226;
 buffer[1158] = 226;
 buffer[1159] = 226;
 buffer[1160] = 225;
 buffer[1161] = 225;
 buffer[1162] = 225;
 buffer[1163] = 225;
 buffer[1164] = 225;
 buffer[1165] = 225;
 buffer[1166] = 224;
 buffer[1167] = 224;
 buffer[1168] = 224;
 buffer[1169] = 224;
 buffer[1170] = 224;
 buffer[1171] = 223;
 buffer[1172] = 223;
 buffer[1173] = 223;
 buffer[1174] = 223;
 buffer[1175] = 223;
 buffer[1176] = 222;
 buffer[1177] = 222;
 buffer[1178] = 222;
 buffer[1179] = 222;
 buffer[1180] = 222;
 buffer[1181] = 221;
 buffer[1182] = 221;
 buffer[1183] = 221;
 buffer[1184] = 221;
 buffer[1185] = 221;
 buffer[1186] = 221;
 buffer[1187] = 220;
 buffer[1188] = 220;
 buffer[1189] = 220;
 buffer[1190] = 220;
 buffer[1191] = 220;
 buffer[1192] = 219;
 buffer[1193] = 219;
 buffer[1194] = 219;
 buffer[1195] = 219;
 buffer[1196] = 219;
 buffer[1197] = 219;
 buffer[1198] = 218;
 buffer[1199] = 218;
 buffer[1200] = 218;
 buffer[1201] = 218;
 buffer[1202] = 218;
 buffer[1203] = 217;
 buffer[1204] = 217;
 buffer[1205] = 217;
 buffer[1206] = 217;
 buffer[1207] = 217;
 buffer[1208] = 217;
 buffer[1209] = 216;
 buffer[1210] = 216;
 buffer[1211] = 216;
 buffer[1212] = 216;
 buffer[1213] = 216;
 buffer[1214] = 215;
 buffer[1215] = 215;
 buffer[1216] = 215;
 buffer[1217] = 215;
 buffer[1218] = 215;
 buffer[1219] = 215;
 buffer[1220] = 214;
 buffer[1221] = 214;
 buffer[1222] = 214;
 buffer[1223] = 214;
 buffer[1224] = 214;
 buffer[1225] = 213;
 buffer[1226] = 213;
 buffer[1227] = 213;
 buffer[1228] = 213;
 buffer[1229] = 213;
 buffer[1230] = 213;
 buffer[1231] = 212;
 buffer[1232] = 212;
 buffer[1233] = 212;
 buffer[1234] = 212;
 buffer[1235] = 212;
 buffer[1236] = 212;
 buffer[1237] = 211;
 buffer[1238] = 211;
 buffer[1239] = 211;
 buffer[1240] = 211;
 buffer[1241] = 211;
 buffer[1242] = 211;
 buffer[1243] = 210;
 buffer[1244] = 210;
 buffer[1245] = 210;
 buffer[1246] = 210;
 buffer[1247] = 210;
 buffer[1248] = 210;
 buffer[1249] = 209;
 buffer[1250] = 209;
 buffer[1251] = 209;
 buffer[1252] = 209;
 buffer[1253] = 209;
 buffer[1254] = 209;
 buffer[1255] = 208;
 buffer[1256] = 208;
 buffer[1257] = 208;
 buffer[1258] = 208;
 buffer[1259] = 208;
 buffer[1260] = 208;
 buffer[1261] = 207;
 buffer[1262] = 207;
 buffer[1263] = 207;
 buffer[1264] = 207;
 buffer[1265] = 207;
 buffer[1266] = 207;
 buffer[1267] = 206;
 buffer[1268] = 206;
 buffer[1269] = 206;
 buffer[1270] = 206;
 buffer[1271] = 206;
 buffer[1272] = 206;
 buffer[1273] = 205;
 buffer[1274] = 205;
 buffer[1275] = 205;
 buffer[1276] = 205;
 buffer[1277] = 205;
 buffer[1278] = 205;
 buffer[1279] = 204;
 buffer[1280] = 204;
 buffer[1281] = 204;
 buffer[1282] = 204;
 buffer[1283] = 204;
 buffer[1284] = 204;
 buffer[1285] = 204;
 buffer[1286] = 203;
 buffer[1287] = 203;
 buffer[1288] = 203;
 buffer[1289] = 203;
 buffer[1290] = 203;
 buffer[1291] = 203;
 buffer[1292] = 202;
 buffer[1293] = 202;
 buffer[1294] = 202;
 buffer[1295] = 202;
 buffer[1296] = 202;
 buffer[1297] = 202;
 buffer[1298] = 201;
 buffer[1299] = 201;
 buffer[1300] = 201;
 buffer[1301] = 201;
 buffer[1302] = 201;
 buffer[1303] = 201;
 buffer[1304] = 201;
 buffer[1305] = 200;
 buffer[1306] = 200;
 buffer[1307] = 200;
 buffer[1308] = 200;
 buffer[1309] = 200;
 buffer[1310] = 200;
 buffer[1311] = 199;
 buffer[1312] = 199;
 buffer[1313] = 199;
 buffer[1314] = 199;
 buffer[1315] = 199;
 buffer[1316] = 199;
 buffer[1317] = 199;
 buffer[1318] = 198;
 buffer[1319] = 198;
 buffer[1320] = 198;
 buffer[1321] = 198;
 buffer[1322] = 198;
 buffer[1323] = 198;
 buffer[1324] = 197;
 buffer[1325] = 197;
 buffer[1326] = 197;
 buffer[1327] = 197;
 buffer[1328] = 197;
 buffer[1329] = 197;
 buffer[1330] = 197;
 buffer[1331] = 196;
 buffer[1332] = 196;
 buffer[1333] = 196;
 buffer[1334] = 196;
 buffer[1335] = 196;
 buffer[1336] = 196;
 buffer[1337] = 196;
 buffer[1338] = 195;
 buffer[1339] = 195;
 buffer[1340] = 195;
 buffer[1341] = 195;
 buffer[1342] = 195;
 buffer[1343] = 195;
 buffer[1344] = 195;
 buffer[1345] = 194;
 buffer[1346] = 194;
 buffer[1347] = 194;
 buffer[1348] = 194;
 buffer[1349] = 194;
 buffer[1350] = 194;
 buffer[1351] = 194;
 buffer[1352] = 193;
 buffer[1353] = 193;
 buffer[1354] = 193;
 buffer[1355] = 193;
 buffer[1356] = 193;
 buffer[1357] = 193;
 buffer[1358] = 193;
 buffer[1359] = 192;
 buffer[1360] = 192;
 buffer[1361] = 192;
 buffer[1362] = 192;
 buffer[1363] = 192;
 buffer[1364] = 192;
 buffer[1365] = 192;
 buffer[1366] = 191;
 buffer[1367] = 191;
 buffer[1368] = 191;
 buffer[1369] = 191;
 buffer[1370] = 191;
 buffer[1371] = 191;
 buffer[1372] = 191;
 buffer[1373] = 190;
 buffer[1374] = 190;
 buffer[1375] = 190;
 buffer[1376] = 190;
 buffer[1377] = 190;
 buffer[1378] = 190;
 buffer[1379] = 190;
 buffer[1380] = 189;
 buffer[1381] = 189;
 buffer[1382] = 189;
 buffer[1383] = 189;
 buffer[1384] = 189;
 buffer[1385] = 189;
 buffer[1386] = 189;
 buffer[1387] = 189;
 buffer[1388] = 188;
 buffer[1389] = 188;
 buffer[1390] = 188;
 buffer[1391] = 188;
 buffer[1392] = 188;
 buffer[1393] = 188;
 buffer[1394] = 188;
 buffer[1395] = 187;
 buffer[1396] = 187;
 buffer[1397] = 187;
 buffer[1398] = 187;
 buffer[1399] = 187;
 buffer[1400] = 187;
 buffer[1401] = 187;
 buffer[1402] = 186;
 buffer[1403] = 186;
 buffer[1404] = 186;
 buffer[1405] = 186;
 buffer[1406] = 186;
 buffer[1407] = 186;
 buffer[1408] = 186;
 buffer[1409] = 186;
 buffer[1410] = 185;
 buffer[1411] = 185;
 buffer[1412] = 185;
 buffer[1413] = 185;
 buffer[1414] = 185;
 buffer[1415] = 185;
 buffer[1416] = 185;
 buffer[1417] = 184;
 buffer[1418] = 184;
 buffer[1419] = 184;
 buffer[1420] = 184;
 buffer[1421] = 184;
 buffer[1422] = 184;
 buffer[1423] = 184;
 buffer[1424] = 184;
 buffer[1425] = 183;
 buffer[1426] = 183;
 buffer[1427] = 183;
 buffer[1428] = 183;
 buffer[1429] = 183;
 buffer[1430] = 183;
 buffer[1431] = 183;
 buffer[1432] = 183;
 buffer[1433] = 182;
 buffer[1434] = 182;
 buffer[1435] = 182;
 buffer[1436] = 182;
 buffer[1437] = 182;
 buffer[1438] = 182;
 buffer[1439] = 182;
 buffer[1440] = 182;
 buffer[1441] = 181;
 buffer[1442] = 181;
 buffer[1443] = 181;
 buffer[1444] = 181;
 buffer[1445] = 181;
 buffer[1446] = 181;
 buffer[1447] = 181;
 buffer[1448] = 181;
 buffer[1449] = 180;
 buffer[1450] = 180;
 buffer[1451] = 180;
 buffer[1452] = 180;
 buffer[1453] = 180;
 buffer[1454] = 180;
 buffer[1455] = 180;
 buffer[1456] = 180;
 buffer[1457] = 179;
 buffer[1458] = 179;
 buffer[1459] = 179;
 buffer[1460] = 179;
 buffer[1461] = 179;
 buffer[1462] = 179;
 buffer[1463] = 179;
 buffer[1464] = 179;
 buffer[1465] = 178;
 buffer[1466] = 178;
 buffer[1467] = 178;
 buffer[1468] = 178;
 buffer[1469] = 178;
 buffer[1470] = 178;
 buffer[1471] = 178;
 buffer[1472] = 178;
 buffer[1473] = 177;
 buffer[1474] = 177;
 buffer[1475] = 177;
 buffer[1476] = 177;
 buffer[1477] = 177;
 buffer[1478] = 177;
 buffer[1479] = 177;
 buffer[1480] = 177;
 buffer[1481] = 177;
 buffer[1482] = 176;
 buffer[1483] = 176;
 buffer[1484] = 176;
 buffer[1485] = 176;
 buffer[1486] = 176;
 buffer[1487] = 176;
 buffer[1488] = 176;
 buffer[1489] = 176;
 buffer[1490] = 175;
 buffer[1491] = 175;
 buffer[1492] = 175;
 buffer[1493] = 175;
 buffer[1494] = 175;
 buffer[1495] = 175;
 buffer[1496] = 175;
 buffer[1497] = 175;
 buffer[1498] = 174;
 buffer[1499] = 174;
 buffer[1500] = 174;
 buffer[1501] = 174;
 buffer[1502] = 174;
 buffer[1503] = 174;
 buffer[1504] = 174;
 buffer[1505] = 174;
 buffer[1506] = 174;
 buffer[1507] = 173;
 buffer[1508] = 173;
 buffer[1509] = 173;
 buffer[1510] = 173;
 buffer[1511] = 173;
 buffer[1512] = 173;
 buffer[1513] = 173;
 buffer[1514] = 173;
 buffer[1515] = 173;
 buffer[1516] = 172;
 buffer[1517] = 172;
 buffer[1518] = 172;
 buffer[1519] = 172;
 buffer[1520] = 172;
 buffer[1521] = 172;
 buffer[1522] = 172;
 buffer[1523] = 172;
 buffer[1524] = 172;
 buffer[1525] = 171;
 buffer[1526] = 171;
 buffer[1527] = 171;
 buffer[1528] = 171;
 buffer[1529] = 171;
 buffer[1530] = 171;
 buffer[1531] = 171;
 buffer[1532] = 171;
 buffer[1533] = 171;
 buffer[1534] = 170;
 buffer[1535] = 170;
 buffer[1536] = 170;
 buffer[1537] = 170;
 buffer[1538] = 170;
 buffer[1539] = 170;
 buffer[1540] = 170;
 buffer[1541] = 170;
 buffer[1542] = 170;
 buffer[1543] = 169;
 buffer[1544] = 169;
 buffer[1545] = 169;
 buffer[1546] = 169;
 buffer[1547] = 169;
 buffer[1548] = 169;
 buffer[1549] = 169;
 buffer[1550] = 169;
 buffer[1551] = 169;
 buffer[1552] = 168;
 buffer[1553] = 168;
 buffer[1554] = 168;
 buffer[1555] = 168;
 buffer[1556] = 168;
 buffer[1557] = 168;
 buffer[1558] = 168;
 buffer[1559] = 168;
 buffer[1560] = 168;
 buffer[1561] = 167;
 buffer[1562] = 167;
 buffer[1563] = 167;
 buffer[1564] = 167;
 buffer[1565] = 167;
 buffer[1566] = 167;
 buffer[1567] = 167;
 buffer[1568] = 167;
 buffer[1569] = 167;
 buffer[1570] = 166;
 buffer[1571] = 166;
 buffer[1572] = 166;
 buffer[1573] = 166;
 buffer[1574] = 166;
 buffer[1575] = 166;
 buffer[1576] = 166;
 buffer[1577] = 166;
 buffer[1578] = 166;
 buffer[1579] = 166;
 buffer[1580] = 165;
 buffer[1581] = 165;
 buffer[1582] = 165;
 buffer[1583] = 165;
 buffer[1584] = 165;
 buffer[1585] = 165;
 buffer[1586] = 165;
 buffer[1587] = 165;
 buffer[1588] = 165;
 buffer[1589] = 164;
 buffer[1590] = 164;
 buffer[1591] = 164;
 buffer[1592] = 164;
 buffer[1593] = 164;
 buffer[1594] = 164;
 buffer[1595] = 164;
 buffer[1596] = 164;
 buffer[1597] = 164;
 buffer[1598] = 164;
 buffer[1599] = 163;
 buffer[1600] = 163;
 buffer[1601] = 163;
 buffer[1602] = 163;
 buffer[1603] = 163;
 buffer[1604] = 163;
 buffer[1605] = 163;
 buffer[1606] = 163;
 buffer[1607] = 163;
 buffer[1608] = 163;
 buffer[1609] = 162;
 buffer[1610] = 162;
 buffer[1611] = 162;
 buffer[1612] = 162;
 buffer[1613] = 162;
 buffer[1614] = 162;
 buffer[1615] = 162;
 buffer[1616] = 162;
 buffer[1617] = 162;
 buffer[1618] = 162;
 buffer[1619] = 161;
 buffer[1620] = 161;
 buffer[1621] = 161;
 buffer[1622] = 161;
 buffer[1623] = 161;
 buffer[1624] = 161;
 buffer[1625] = 161;
 buffer[1626] = 161;
 buffer[1627] = 161;
 buffer[1628] = 161;
 buffer[1629] = 160;
 buffer[1630] = 160;
 buffer[1631] = 160;
 buffer[1632] = 160;
 buffer[1633] = 160;
 buffer[1634] = 160;
 buffer[1635] = 160;
 buffer[1636] = 160;
 buffer[1637] = 160;
 buffer[1638] = 160;
 buffer[1639] = 159;
 buffer[1640] = 159;
 buffer[1641] = 159;
 buffer[1642] = 159;
 buffer[1643] = 159;
 buffer[1644] = 159;
 buffer[1645] = 159;
 buffer[1646] = 159;
 buffer[1647] = 159;
 buffer[1648] = 159;
 buffer[1649] = 158;
 buffer[1650] = 158;
 buffer[1651] = 158;
 buffer[1652] = 158;
 buffer[1653] = 158;
 buffer[1654] = 158;
 buffer[1655] = 158;
 buffer[1656] = 158;
 buffer[1657] = 158;
 buffer[1658] = 158;
 buffer[1659] = 158;
 buffer[1660] = 157;
 buffer[1661] = 157;
 buffer[1662] = 157;
 buffer[1663] = 157;
 buffer[1664] = 157;
 buffer[1665] = 157;
 buffer[1666] = 157;
 buffer[1667] = 157;
 buffer[1668] = 157;
 buffer[1669] = 157;
 buffer[1670] = 156;
 buffer[1671] = 156;
 buffer[1672] = 156;
 buffer[1673] = 156;
 buffer[1674] = 156;
 buffer[1675] = 156;
 buffer[1676] = 156;
 buffer[1677] = 156;
 buffer[1678] = 156;
 buffer[1679] = 156;
 buffer[1680] = 156;
 buffer[1681] = 155;
 buffer[1682] = 155;
 buffer[1683] = 155;
 buffer[1684] = 155;
 buffer[1685] = 155;
 buffer[1686] = 155;
 buffer[1687] = 155;
 buffer[1688] = 155;
 buffer[1689] = 155;
 buffer[1690] = 155;
 buffer[1691] = 155;
 buffer[1692] = 154;
 buffer[1693] = 154;
 buffer[1694] = 154;
 buffer[1695] = 154;
 buffer[1696] = 154;
 buffer[1697] = 154;
 buffer[1698] = 154;
 buffer[1699] = 154;
 buffer[1700] = 154;
 buffer[1701] = 154;
 buffer[1702] = 154;
 buffer[1703] = 153;
 buffer[1704] = 153;
 buffer[1705] = 153;
 buffer[1706] = 153;
 buffer[1707] = 153;
 buffer[1708] = 153;
 buffer[1709] = 153;
 buffer[1710] = 153;
 buffer[1711] = 153;
 buffer[1712] = 153;
 buffer[1713] = 153;
 buffer[1714] = 152;
 buffer[1715] = 152;
 buffer[1716] = 152;
 buffer[1717] = 152;
 buffer[1718] = 152;
 buffer[1719] = 152;
 buffer[1720] = 152;
 buffer[1721] = 152;
 buffer[1722] = 152;
 buffer[1723] = 152;
 buffer[1724] = 152;
 buffer[1725] = 151;
 buffer[1726] = 151;
 buffer[1727] = 151;
 buffer[1728] = 151;
 buffer[1729] = 151;
 buffer[1730] = 151;
 buffer[1731] = 151;
 buffer[1732] = 151;
 buffer[1733] = 151;
 buffer[1734] = 151;
 buffer[1735] = 151;
 buffer[1736] = 151;
 buffer[1737] = 150;
 buffer[1738] = 150;
 buffer[1739] = 150;
 buffer[1740] = 150;
 buffer[1741] = 150;
 buffer[1742] = 150;
 buffer[1743] = 150;
 buffer[1744] = 150;
 buffer[1745] = 150;
 buffer[1746] = 150;
 buffer[1747] = 150;
 buffer[1748] = 149;
 buffer[1749] = 149;
 buffer[1750] = 149;
 buffer[1751] = 149;
 buffer[1752] = 149;
 buffer[1753] = 149;
 buffer[1754] = 149;
 buffer[1755] = 149;
 buffer[1756] = 149;
 buffer[1757] = 149;
 buffer[1758] = 149;
 buffer[1759] = 149;
 buffer[1760] = 148;
 buffer[1761] = 148;
 buffer[1762] = 148;
 buffer[1763] = 148;
 buffer[1764] = 148;
 buffer[1765] = 148;
 buffer[1766] = 148;
 buffer[1767] = 148;
 buffer[1768] = 148;
 buffer[1769] = 148;
 buffer[1770] = 148;
 buffer[1771] = 148;
 buffer[1772] = 147;
 buffer[1773] = 147;
 buffer[1774] = 147;
 buffer[1775] = 147;
 buffer[1776] = 147;
 buffer[1777] = 147;
 buffer[1778] = 147;
 buffer[1779] = 147;
 buffer[1780] = 147;
 buffer[1781] = 147;
 buffer[1782] = 147;
 buffer[1783] = 147;
 buffer[1784] = 146;
 buffer[1785] = 146;
 buffer[1786] = 146;
 buffer[1787] = 146;
 buffer[1788] = 146;
 buffer[1789] = 146;
 buffer[1790] = 146;
 buffer[1791] = 146;
 buffer[1792] = 146;
 buffer[1793] = 146;
 buffer[1794] = 146;
 buffer[1795] = 146;
 buffer[1796] = 145;
 buffer[1797] = 145;
 buffer[1798] = 145;
 buffer[1799] = 145;
 buffer[1800] = 145;
 buffer[1801] = 145;
 buffer[1802] = 145;
 buffer[1803] = 145;
 buffer[1804] = 145;
 buffer[1805] = 145;
 buffer[1806] = 145;
 buffer[1807] = 145;
 buffer[1808] = 144;
 buffer[1809] = 144;
 buffer[1810] = 144;
 buffer[1811] = 144;
 buffer[1812] = 144;
 buffer[1813] = 144;
 buffer[1814] = 144;
 buffer[1815] = 144;
 buffer[1816] = 144;
 buffer[1817] = 144;
 buffer[1818] = 144;
 buffer[1819] = 144;
 buffer[1820] = 144;
 buffer[1821] = 143;
 buffer[1822] = 143;
 buffer[1823] = 143;
 buffer[1824] = 143;
 buffer[1825] = 143;
 buffer[1826] = 143;
 buffer[1827] = 143;
 buffer[1828] = 143;
 buffer[1829] = 143;
 buffer[1830] = 143;
 buffer[1831] = 143;
 buffer[1832] = 143;
 buffer[1833] = 143;
 buffer[1834] = 142;
 buffer[1835] = 142;
 buffer[1836] = 142;
 buffer[1837] = 142;
 buffer[1838] = 142;
 buffer[1839] = 142;
 buffer[1840] = 142;
 buffer[1841] = 142;
 buffer[1842] = 142;
 buffer[1843] = 142;
 buffer[1844] = 142;
 buffer[1845] = 142;
 buffer[1846] = 142;
 buffer[1847] = 141;
 buffer[1848] = 141;
 buffer[1849] = 141;
 buffer[1850] = 141;
 buffer[1851] = 141;
 buffer[1852] = 141;
 buffer[1853] = 141;
 buffer[1854] = 141;
 buffer[1855] = 141;
 buffer[1856] = 141;
 buffer[1857] = 141;
 buffer[1858] = 141;
 buffer[1859] = 141;
 buffer[1860] = 140;
 buffer[1861] = 140;
 buffer[1862] = 140;
 buffer[1863] = 140;
 buffer[1864] = 140;
 buffer[1865] = 140;
 buffer[1866] = 140;
 buffer[1867] = 140;
 buffer[1868] = 140;
 buffer[1869] = 140;
 buffer[1870] = 140;
 buffer[1871] = 140;
 buffer[1872] = 140;
 buffer[1873] = 139;
 buffer[1874] = 139;
 buffer[1875] = 139;
 buffer[1876] = 139;
 buffer[1877] = 139;
 buffer[1878] = 139;
 buffer[1879] = 139;
 buffer[1880] = 139;
 buffer[1881] = 139;
 buffer[1882] = 139;
 buffer[1883] = 139;
 buffer[1884] = 139;
 buffer[1885] = 139;
 buffer[1886] = 138;
 buffer[1887] = 138;
 buffer[1888] = 138;
 buffer[1889] = 138;
 buffer[1890] = 138;
 buffer[1891] = 138;
 buffer[1892] = 138;
 buffer[1893] = 138;
 buffer[1894] = 138;
 buffer[1895] = 138;
 buffer[1896] = 138;
 buffer[1897] = 138;
 buffer[1898] = 138;
 buffer[1899] = 138;
 buffer[1900] = 137;
 buffer[1901] = 137;
 buffer[1902] = 137;
 buffer[1903] = 137;
 buffer[1904] = 137;
 buffer[1905] = 137;
 buffer[1906] = 137;
 buffer[1907] = 137;
 buffer[1908] = 137;
 buffer[1909] = 137;
 buffer[1910] = 137;
 buffer[1911] = 137;
 buffer[1912] = 137;
 buffer[1913] = 137;
 buffer[1914] = 136;
 buffer[1915] = 136;
 buffer[1916] = 136;
 buffer[1917] = 136;
 buffer[1918] = 136;
 buffer[1919] = 136;
 buffer[1920] = 136;
 buffer[1921] = 136;
 buffer[1922] = 136;
 buffer[1923] = 136;
 buffer[1924] = 136;
 buffer[1925] = 136;
 buffer[1926] = 136;
 buffer[1927] = 136;
 buffer[1928] = 135;
 buffer[1929] = 135;
 buffer[1930] = 135;
 buffer[1931] = 135;
 buffer[1932] = 135;
 buffer[1933] = 135;
 buffer[1934] = 135;
 buffer[1935] = 135;
 buffer[1936] = 135;
 buffer[1937] = 135;
 buffer[1938] = 135;
 buffer[1939] = 135;
 buffer[1940] = 135;
 buffer[1941] = 135;
 buffer[1942] = 134;
 buffer[1943] = 134;
 buffer[1944] = 134;
 buffer[1945] = 134;
 buffer[1946] = 134;
 buffer[1947] = 134;
 buffer[1948] = 134;
 buffer[1949] = 134;
 buffer[1950] = 134;
 buffer[1951] = 134;
 buffer[1952] = 134;
 buffer[1953] = 134;
 buffer[1954] = 134;
 buffer[1955] = 134;
 buffer[1956] = 134;
 buffer[1957] = 133;
 buffer[1958] = 133;
 buffer[1959] = 133;
 buffer[1960] = 133;
 buffer[1961] = 133;
 buffer[1962] = 133;
 buffer[1963] = 133;
 buffer[1964] = 133;
 buffer[1965] = 133;
 buffer[1966] = 133;
 buffer[1967] = 133;
 buffer[1968] = 133;
 buffer[1969] = 133;
 buffer[1970] = 133;
 buffer[1971] = 133;
 buffer[1972] = 132;
 buffer[1973] = 132;
 buffer[1974] = 132;
 buffer[1975] = 132;
 buffer[1976] = 132;
 buffer[1977] = 132;
 buffer[1978] = 132;
 buffer[1979] = 132;
 buffer[1980] = 132;
 buffer[1981] = 132;
 buffer[1982] = 132;
 buffer[1983] = 132;
 buffer[1984] = 132;
 buffer[1985] = 132;
 buffer[1986] = 131;
 buffer[1987] = 131;
 buffer[1988] = 131;
 buffer[1989] = 131;
 buffer[1990] = 131;
 buffer[1991] = 131;
 buffer[1992] = 131;
 buffer[1993] = 131;
 buffer[1994] = 131;
 buffer[1995] = 131;
 buffer[1996] = 131;
 buffer[1997] = 131;
 buffer[1998] = 131;
 buffer[1999] = 131;
 buffer[2000] = 131;
 buffer[2001] = 131;
 buffer[2002] = 130;
 buffer[2003] = 130;
 buffer[2004] = 130;
 buffer[2005] = 130;
 buffer[2006] = 130;
 buffer[2007] = 130;
 buffer[2008] = 130;
 buffer[2009] = 130;
 buffer[2010] = 130;
 buffer[2011] = 130;
 buffer[2012] = 130;
 buffer[2013] = 130;
 buffer[2014] = 130;
 buffer[2015] = 130;
 buffer[2016] = 130;
 buffer[2017] = 129;
 buffer[2018] = 129;
 buffer[2019] = 129;
 buffer[2020] = 129;
 buffer[2021] = 129;
 buffer[2022] = 129;
 buffer[2023] = 129;
 buffer[2024] = 129;
 buffer[2025] = 129;
 buffer[2026] = 129;
 buffer[2027] = 129;
 buffer[2028] = 129;
 buffer[2029] = 129;
 buffer[2030] = 129;
 buffer[2031] = 129;
 buffer[2032] = 129;
 buffer[2033] = 128;
 buffer[2034] = 128;
 buffer[2035] = 128;
 buffer[2036] = 128;
 buffer[2037] = 128;
 buffer[2038] = 128;
 buffer[2039] = 128;
 buffer[2040] = 128;
 buffer[2041] = 128;
 buffer[2042] = 128;
 buffer[2043] = 128;
 buffer[2044] = 128;
 buffer[2045] = 128;
 buffer[2046] = 128;
 buffer[2047] = 128;
end

endmodule

// SL 2019, MIT license
module M_frame_display__mem_invB(
input                  [1-1:0] in_wenable,
input       [18-1:0]    in_wdata,
input                  [11-1:0]    in_addr,
output reg  [18-1:0]    out_rdata,
input                                        clock
);
  (* no_rw_check *) reg  [18-1:0] buffer[2048-1:0];
`ifdef SIMULATION
  // in simulation we use a different code that matches yosys output with
  // no_rw_check enabled (which we use to preserve compact LUT designs)
  always @(posedge clock) begin
    if (in_wenable) begin
      buffer[in_addr] <= in_wdata;
      out_rdata       <= in_wdata;
    end else begin
      out_rdata       <= buffer[in_addr];
    end
  end
`else
  always @(posedge clock) begin
    if (in_wenable) begin
      buffer[in_addr] <= in_wdata;
    end
    out_rdata <= buffer[in_addr];
  end
`endif
initial begin
 buffer[0] = 131071;
 buffer[1] = 131071;
 buffer[2] = 131071;
 buffer[3] = 87381;
 buffer[4] = 65536;
 buffer[5] = 52428;
 buffer[6] = 43690;
 buffer[7] = 37449;
 buffer[8] = 32768;
 buffer[9] = 29127;
 buffer[10] = 26214;
 buffer[11] = 23831;
 buffer[12] = 21845;
 buffer[13] = 20164;
 buffer[14] = 18724;
 buffer[15] = 17476;
 buffer[16] = 16384;
 buffer[17] = 15420;
 buffer[18] = 14563;
 buffer[19] = 13797;
 buffer[20] = 13107;
 buffer[21] = 12483;
 buffer[22] = 11915;
 buffer[23] = 11397;
 buffer[24] = 10922;
 buffer[25] = 10485;
 buffer[26] = 10082;
 buffer[27] = 9709;
 buffer[28] = 9362;
 buffer[29] = 9039;
 buffer[30] = 8738;
 buffer[31] = 8456;
 buffer[32] = 8192;
 buffer[33] = 7943;
 buffer[34] = 7710;
 buffer[35] = 7489;
 buffer[36] = 7281;
 buffer[37] = 7084;
 buffer[38] = 6898;
 buffer[39] = 6721;
 buffer[40] = 6553;
 buffer[41] = 6393;
 buffer[42] = 6241;
 buffer[43] = 6096;
 buffer[44] = 5957;
 buffer[45] = 5825;
 buffer[46] = 5698;
 buffer[47] = 5577;
 buffer[48] = 5461;
 buffer[49] = 5349;
 buffer[50] = 5242;
 buffer[51] = 5140;
 buffer[52] = 5041;
 buffer[53] = 4946;
 buffer[54] = 4854;
 buffer[55] = 4766;
 buffer[56] = 4681;
 buffer[57] = 4599;
 buffer[58] = 4519;
 buffer[59] = 4443;
 buffer[60] = 4369;
 buffer[61] = 4297;
 buffer[62] = 4228;
 buffer[63] = 4161;
 buffer[64] = 4096;
 buffer[65] = 4032;
 buffer[66] = 3971;
 buffer[67] = 3912;
 buffer[68] = 3855;
 buffer[69] = 3799;
 buffer[70] = 3744;
 buffer[71] = 3692;
 buffer[72] = 3640;
 buffer[73] = 3591;
 buffer[74] = 3542;
 buffer[75] = 3495;
 buffer[76] = 3449;
 buffer[77] = 3404;
 buffer[78] = 3360;
 buffer[79] = 3318;
 buffer[80] = 3276;
 buffer[81] = 3236;
 buffer[82] = 3196;
 buffer[83] = 3158;
 buffer[84] = 3120;
 buffer[85] = 3084;
 buffer[86] = 3048;
 buffer[87] = 3013;
 buffer[88] = 2978;
 buffer[89] = 2945;
 buffer[90] = 2912;
 buffer[91] = 2880;
 buffer[92] = 2849;
 buffer[93] = 2818;
 buffer[94] = 2788;
 buffer[95] = 2759;
 buffer[96] = 2730;
 buffer[97] = 2702;
 buffer[98] = 2674;
 buffer[99] = 2647;
 buffer[100] = 2621;
 buffer[101] = 2595;
 buffer[102] = 2570;
 buffer[103] = 2545;
 buffer[104] = 2520;
 buffer[105] = 2496;
 buffer[106] = 2473;
 buffer[107] = 2449;
 buffer[108] = 2427;
 buffer[109] = 2404;
 buffer[110] = 2383;
 buffer[111] = 2361;
 buffer[112] = 2340;
 buffer[113] = 2319;
 buffer[114] = 2299;
 buffer[115] = 2279;
 buffer[116] = 2259;
 buffer[117] = 2240;
 buffer[118] = 2221;
 buffer[119] = 2202;
 buffer[120] = 2184;
 buffer[121] = 2166;
 buffer[122] = 2148;
 buffer[123] = 2131;
 buffer[124] = 2114;
 buffer[125] = 2097;
 buffer[126] = 2080;
 buffer[127] = 2064;
 buffer[128] = 2048;
 buffer[129] = 2032;
 buffer[130] = 2016;
 buffer[131] = 2001;
 buffer[132] = 1985;
 buffer[133] = 1971;
 buffer[134] = 1956;
 buffer[135] = 1941;
 buffer[136] = 1927;
 buffer[137] = 1913;
 buffer[138] = 1899;
 buffer[139] = 1885;
 buffer[140] = 1872;
 buffer[141] = 1859;
 buffer[142] = 1846;
 buffer[143] = 1833;
 buffer[144] = 1820;
 buffer[145] = 1807;
 buffer[146] = 1795;
 buffer[147] = 1783;
 buffer[148] = 1771;
 buffer[149] = 1759;
 buffer[150] = 1747;
 buffer[151] = 1736;
 buffer[152] = 1724;
 buffer[153] = 1713;
 buffer[154] = 1702;
 buffer[155] = 1691;
 buffer[156] = 1680;
 buffer[157] = 1669;
 buffer[158] = 1659;
 buffer[159] = 1648;
 buffer[160] = 1638;
 buffer[161] = 1628;
 buffer[162] = 1618;
 buffer[163] = 1608;
 buffer[164] = 1598;
 buffer[165] = 1588;
 buffer[166] = 1579;
 buffer[167] = 1569;
 buffer[168] = 1560;
 buffer[169] = 1551;
 buffer[170] = 1542;
 buffer[171] = 1533;
 buffer[172] = 1524;
 buffer[173] = 1515;
 buffer[174] = 1506;
 buffer[175] = 1497;
 buffer[176] = 1489;
 buffer[177] = 1481;
 buffer[178] = 1472;
 buffer[179] = 1464;
 buffer[180] = 1456;
 buffer[181] = 1448;
 buffer[182] = 1440;
 buffer[183] = 1432;
 buffer[184] = 1424;
 buffer[185] = 1416;
 buffer[186] = 1409;
 buffer[187] = 1401;
 buffer[188] = 1394;
 buffer[189] = 1387;
 buffer[190] = 1379;
 buffer[191] = 1372;
 buffer[192] = 1365;
 buffer[193] = 1358;
 buffer[194] = 1351;
 buffer[195] = 1344;
 buffer[196] = 1337;
 buffer[197] = 1330;
 buffer[198] = 1323;
 buffer[199] = 1317;
 buffer[200] = 1310;
 buffer[201] = 1304;
 buffer[202] = 1297;
 buffer[203] = 1291;
 buffer[204] = 1285;
 buffer[205] = 1278;
 buffer[206] = 1272;
 buffer[207] = 1266;
 buffer[208] = 1260;
 buffer[209] = 1254;
 buffer[210] = 1248;
 buffer[211] = 1242;
 buffer[212] = 1236;
 buffer[213] = 1230;
 buffer[214] = 1224;
 buffer[215] = 1219;
 buffer[216] = 1213;
 buffer[217] = 1208;
 buffer[218] = 1202;
 buffer[219] = 1197;
 buffer[220] = 1191;
 buffer[221] = 1186;
 buffer[222] = 1180;
 buffer[223] = 1175;
 buffer[224] = 1170;
 buffer[225] = 1165;
 buffer[226] = 1159;
 buffer[227] = 1154;
 buffer[228] = 1149;
 buffer[229] = 1144;
 buffer[230] = 1139;
 buffer[231] = 1134;
 buffer[232] = 1129;
 buffer[233] = 1125;
 buffer[234] = 1120;
 buffer[235] = 1115;
 buffer[236] = 1110;
 buffer[237] = 1106;
 buffer[238] = 1101;
 buffer[239] = 1096;
 buffer[240] = 1092;
 buffer[241] = 1087;
 buffer[242] = 1083;
 buffer[243] = 1078;
 buffer[244] = 1074;
 buffer[245] = 1069;
 buffer[246] = 1065;
 buffer[247] = 1061;
 buffer[248] = 1057;
 buffer[249] = 1052;
 buffer[250] = 1048;
 buffer[251] = 1044;
 buffer[252] = 1040;
 buffer[253] = 1036;
 buffer[254] = 1032;
 buffer[255] = 1028;
 buffer[256] = 1024;
 buffer[257] = 1020;
 buffer[258] = 1016;
 buffer[259] = 1012;
 buffer[260] = 1008;
 buffer[261] = 1004;
 buffer[262] = 1000;
 buffer[263] = 996;
 buffer[264] = 992;
 buffer[265] = 989;
 buffer[266] = 985;
 buffer[267] = 981;
 buffer[268] = 978;
 buffer[269] = 974;
 buffer[270] = 970;
 buffer[271] = 967;
 buffer[272] = 963;
 buffer[273] = 960;
 buffer[274] = 956;
 buffer[275] = 953;
 buffer[276] = 949;
 buffer[277] = 946;
 buffer[278] = 942;
 buffer[279] = 939;
 buffer[280] = 936;
 buffer[281] = 932;
 buffer[282] = 929;
 buffer[283] = 926;
 buffer[284] = 923;
 buffer[285] = 919;
 buffer[286] = 916;
 buffer[287] = 913;
 buffer[288] = 910;
 buffer[289] = 907;
 buffer[290] = 903;
 buffer[291] = 900;
 buffer[292] = 897;
 buffer[293] = 894;
 buffer[294] = 891;
 buffer[295] = 888;
 buffer[296] = 885;
 buffer[297] = 882;
 buffer[298] = 879;
 buffer[299] = 876;
 buffer[300] = 873;
 buffer[301] = 870;
 buffer[302] = 868;
 buffer[303] = 865;
 buffer[304] = 862;
 buffer[305] = 859;
 buffer[306] = 856;
 buffer[307] = 853;
 buffer[308] = 851;
 buffer[309] = 848;
 buffer[310] = 845;
 buffer[311] = 842;
 buffer[312] = 840;
 buffer[313] = 837;
 buffer[314] = 834;
 buffer[315] = 832;
 buffer[316] = 829;
 buffer[317] = 826;
 buffer[318] = 824;
 buffer[319] = 821;
 buffer[320] = 819;
 buffer[321] = 816;
 buffer[322] = 814;
 buffer[323] = 811;
 buffer[324] = 809;
 buffer[325] = 806;
 buffer[326] = 804;
 buffer[327] = 801;
 buffer[328] = 799;
 buffer[329] = 796;
 buffer[330] = 794;
 buffer[331] = 791;
 buffer[332] = 789;
 buffer[333] = 787;
 buffer[334] = 784;
 buffer[335] = 782;
 buffer[336] = 780;
 buffer[337] = 777;
 buffer[338] = 775;
 buffer[339] = 773;
 buffer[340] = 771;
 buffer[341] = 768;
 buffer[342] = 766;
 buffer[343] = 764;
 buffer[344] = 762;
 buffer[345] = 759;
 buffer[346] = 757;
 buffer[347] = 755;
 buffer[348] = 753;
 buffer[349] = 751;
 buffer[350] = 748;
 buffer[351] = 746;
 buffer[352] = 744;
 buffer[353] = 742;
 buffer[354] = 740;
 buffer[355] = 738;
 buffer[356] = 736;
 buffer[357] = 734;
 buffer[358] = 732;
 buffer[359] = 730;
 buffer[360] = 728;
 buffer[361] = 726;
 buffer[362] = 724;
 buffer[363] = 722;
 buffer[364] = 720;
 buffer[365] = 718;
 buffer[366] = 716;
 buffer[367] = 714;
 buffer[368] = 712;
 buffer[369] = 710;
 buffer[370] = 708;
 buffer[371] = 706;
 buffer[372] = 704;
 buffer[373] = 702;
 buffer[374] = 700;
 buffer[375] = 699;
 buffer[376] = 697;
 buffer[377] = 695;
 buffer[378] = 693;
 buffer[379] = 691;
 buffer[380] = 689;
 buffer[381] = 688;
 buffer[382] = 686;
 buffer[383] = 684;
 buffer[384] = 682;
 buffer[385] = 680;
 buffer[386] = 679;
 buffer[387] = 677;
 buffer[388] = 675;
 buffer[389] = 673;
 buffer[390] = 672;
 buffer[391] = 670;
 buffer[392] = 668;
 buffer[393] = 667;
 buffer[394] = 665;
 buffer[395] = 663;
 buffer[396] = 661;
 buffer[397] = 660;
 buffer[398] = 658;
 buffer[399] = 657;
 buffer[400] = 655;
 buffer[401] = 653;
 buffer[402] = 652;
 buffer[403] = 650;
 buffer[404] = 648;
 buffer[405] = 647;
 buffer[406] = 645;
 buffer[407] = 644;
 buffer[408] = 642;
 buffer[409] = 640;
 buffer[410] = 639;
 buffer[411] = 637;
 buffer[412] = 636;
 buffer[413] = 634;
 buffer[414] = 633;
 buffer[415] = 631;
 buffer[416] = 630;
 buffer[417] = 628;
 buffer[418] = 627;
 buffer[419] = 625;
 buffer[420] = 624;
 buffer[421] = 622;
 buffer[422] = 621;
 buffer[423] = 619;
 buffer[424] = 618;
 buffer[425] = 616;
 buffer[426] = 615;
 buffer[427] = 613;
 buffer[428] = 612;
 buffer[429] = 611;
 buffer[430] = 609;
 buffer[431] = 608;
 buffer[432] = 606;
 buffer[433] = 605;
 buffer[434] = 604;
 buffer[435] = 602;
 buffer[436] = 601;
 buffer[437] = 599;
 buffer[438] = 598;
 buffer[439] = 597;
 buffer[440] = 595;
 buffer[441] = 594;
 buffer[442] = 593;
 buffer[443] = 591;
 buffer[444] = 590;
 buffer[445] = 589;
 buffer[446] = 587;
 buffer[447] = 586;
 buffer[448] = 585;
 buffer[449] = 583;
 buffer[450] = 582;
 buffer[451] = 581;
 buffer[452] = 579;
 buffer[453] = 578;
 buffer[454] = 577;
 buffer[455] = 576;
 buffer[456] = 574;
 buffer[457] = 573;
 buffer[458] = 572;
 buffer[459] = 571;
 buffer[460] = 569;
 buffer[461] = 568;
 buffer[462] = 567;
 buffer[463] = 566;
 buffer[464] = 564;
 buffer[465] = 563;
 buffer[466] = 562;
 buffer[467] = 561;
 buffer[468] = 560;
 buffer[469] = 558;
 buffer[470] = 557;
 buffer[471] = 556;
 buffer[472] = 555;
 buffer[473] = 554;
 buffer[474] = 553;
 buffer[475] = 551;
 buffer[476] = 550;
 buffer[477] = 549;
 buffer[478] = 548;
 buffer[479] = 547;
 buffer[480] = 546;
 buffer[481] = 544;
 buffer[482] = 543;
 buffer[483] = 542;
 buffer[484] = 541;
 buffer[485] = 540;
 buffer[486] = 539;
 buffer[487] = 538;
 buffer[488] = 537;
 buffer[489] = 536;
 buffer[490] = 534;
 buffer[491] = 533;
 buffer[492] = 532;
 buffer[493] = 531;
 buffer[494] = 530;
 buffer[495] = 529;
 buffer[496] = 528;
 buffer[497] = 527;
 buffer[498] = 526;
 buffer[499] = 525;
 buffer[500] = 524;
 buffer[501] = 523;
 buffer[502] = 522;
 buffer[503] = 521;
 buffer[504] = 520;
 buffer[505] = 519;
 buffer[506] = 518;
 buffer[507] = 517;
 buffer[508] = 516;
 buffer[509] = 515;
 buffer[510] = 514;
 buffer[511] = 513;
 buffer[512] = 512;
 buffer[513] = 511;
 buffer[514] = 510;
 buffer[515] = 509;
 buffer[516] = 508;
 buffer[517] = 507;
 buffer[518] = 506;
 buffer[519] = 505;
 buffer[520] = 504;
 buffer[521] = 503;
 buffer[522] = 502;
 buffer[523] = 501;
 buffer[524] = 500;
 buffer[525] = 499;
 buffer[526] = 498;
 buffer[527] = 497;
 buffer[528] = 496;
 buffer[529] = 495;
 buffer[530] = 494;
 buffer[531] = 493;
 buffer[532] = 492;
 buffer[533] = 491;
 buffer[534] = 490;
 buffer[535] = 489;
 buffer[536] = 489;
 buffer[537] = 488;
 buffer[538] = 487;
 buffer[539] = 486;
 buffer[540] = 485;
 buffer[541] = 484;
 buffer[542] = 483;
 buffer[543] = 482;
 buffer[544] = 481;
 buffer[545] = 480;
 buffer[546] = 480;
 buffer[547] = 479;
 buffer[548] = 478;
 buffer[549] = 477;
 buffer[550] = 476;
 buffer[551] = 475;
 buffer[552] = 474;
 buffer[553] = 474;
 buffer[554] = 473;
 buffer[555] = 472;
 buffer[556] = 471;
 buffer[557] = 470;
 buffer[558] = 469;
 buffer[559] = 468;
 buffer[560] = 468;
 buffer[561] = 467;
 buffer[562] = 466;
 buffer[563] = 465;
 buffer[564] = 464;
 buffer[565] = 463;
 buffer[566] = 463;
 buffer[567] = 462;
 buffer[568] = 461;
 buffer[569] = 460;
 buffer[570] = 459;
 buffer[571] = 459;
 buffer[572] = 458;
 buffer[573] = 457;
 buffer[574] = 456;
 buffer[575] = 455;
 buffer[576] = 455;
 buffer[577] = 454;
 buffer[578] = 453;
 buffer[579] = 452;
 buffer[580] = 451;
 buffer[581] = 451;
 buffer[582] = 450;
 buffer[583] = 449;
 buffer[584] = 448;
 buffer[585] = 448;
 buffer[586] = 447;
 buffer[587] = 446;
 buffer[588] = 445;
 buffer[589] = 445;
 buffer[590] = 444;
 buffer[591] = 443;
 buffer[592] = 442;
 buffer[593] = 442;
 buffer[594] = 441;
 buffer[595] = 440;
 buffer[596] = 439;
 buffer[597] = 439;
 buffer[598] = 438;
 buffer[599] = 437;
 buffer[600] = 436;
 buffer[601] = 436;
 buffer[602] = 435;
 buffer[603] = 434;
 buffer[604] = 434;
 buffer[605] = 433;
 buffer[606] = 432;
 buffer[607] = 431;
 buffer[608] = 431;
 buffer[609] = 430;
 buffer[610] = 429;
 buffer[611] = 429;
 buffer[612] = 428;
 buffer[613] = 427;
 buffer[614] = 426;
 buffer[615] = 426;
 buffer[616] = 425;
 buffer[617] = 424;
 buffer[618] = 424;
 buffer[619] = 423;
 buffer[620] = 422;
 buffer[621] = 422;
 buffer[622] = 421;
 buffer[623] = 420;
 buffer[624] = 420;
 buffer[625] = 419;
 buffer[626] = 418;
 buffer[627] = 418;
 buffer[628] = 417;
 buffer[629] = 416;
 buffer[630] = 416;
 buffer[631] = 415;
 buffer[632] = 414;
 buffer[633] = 414;
 buffer[634] = 413;
 buffer[635] = 412;
 buffer[636] = 412;
 buffer[637] = 411;
 buffer[638] = 410;
 buffer[639] = 410;
 buffer[640] = 409;
 buffer[641] = 408;
 buffer[642] = 408;
 buffer[643] = 407;
 buffer[644] = 407;
 buffer[645] = 406;
 buffer[646] = 405;
 buffer[647] = 405;
 buffer[648] = 404;
 buffer[649] = 403;
 buffer[650] = 403;
 buffer[651] = 402;
 buffer[652] = 402;
 buffer[653] = 401;
 buffer[654] = 400;
 buffer[655] = 400;
 buffer[656] = 399;
 buffer[657] = 399;
 buffer[658] = 398;
 buffer[659] = 397;
 buffer[660] = 397;
 buffer[661] = 396;
 buffer[662] = 395;
 buffer[663] = 395;
 buffer[664] = 394;
 buffer[665] = 394;
 buffer[666] = 393;
 buffer[667] = 393;
 buffer[668] = 392;
 buffer[669] = 391;
 buffer[670] = 391;
 buffer[671] = 390;
 buffer[672] = 390;
 buffer[673] = 389;
 buffer[674] = 388;
 buffer[675] = 388;
 buffer[676] = 387;
 buffer[677] = 387;
 buffer[678] = 386;
 buffer[679] = 386;
 buffer[680] = 385;
 buffer[681] = 384;
 buffer[682] = 384;
 buffer[683] = 383;
 buffer[684] = 383;
 buffer[685] = 382;
 buffer[686] = 382;
 buffer[687] = 381;
 buffer[688] = 381;
 buffer[689] = 380;
 buffer[690] = 379;
 buffer[691] = 379;
 buffer[692] = 378;
 buffer[693] = 378;
 buffer[694] = 377;
 buffer[695] = 377;
 buffer[696] = 376;
 buffer[697] = 376;
 buffer[698] = 375;
 buffer[699] = 375;
 buffer[700] = 374;
 buffer[701] = 373;
 buffer[702] = 373;
 buffer[703] = 372;
 buffer[704] = 372;
 buffer[705] = 371;
 buffer[706] = 371;
 buffer[707] = 370;
 buffer[708] = 370;
 buffer[709] = 369;
 buffer[710] = 369;
 buffer[711] = 368;
 buffer[712] = 368;
 buffer[713] = 367;
 buffer[714] = 367;
 buffer[715] = 366;
 buffer[716] = 366;
 buffer[717] = 365;
 buffer[718] = 365;
 buffer[719] = 364;
 buffer[720] = 364;
 buffer[721] = 363;
 buffer[722] = 363;
 buffer[723] = 362;
 buffer[724] = 362;
 buffer[725] = 361;
 buffer[726] = 361;
 buffer[727] = 360;
 buffer[728] = 360;
 buffer[729] = 359;
 buffer[730] = 359;
 buffer[731] = 358;
 buffer[732] = 358;
 buffer[733] = 357;
 buffer[734] = 357;
 buffer[735] = 356;
 buffer[736] = 356;
 buffer[737] = 355;
 buffer[738] = 355;
 buffer[739] = 354;
 buffer[740] = 354;
 buffer[741] = 353;
 buffer[742] = 353;
 buffer[743] = 352;
 buffer[744] = 352;
 buffer[745] = 351;
 buffer[746] = 351;
 buffer[747] = 350;
 buffer[748] = 350;
 buffer[749] = 349;
 buffer[750] = 349;
 buffer[751] = 349;
 buffer[752] = 348;
 buffer[753] = 348;
 buffer[754] = 347;
 buffer[755] = 347;
 buffer[756] = 346;
 buffer[757] = 346;
 buffer[758] = 345;
 buffer[759] = 345;
 buffer[760] = 344;
 buffer[761] = 344;
 buffer[762] = 344;
 buffer[763] = 343;
 buffer[764] = 343;
 buffer[765] = 342;
 buffer[766] = 342;
 buffer[767] = 341;
 buffer[768] = 341;
 buffer[769] = 340;
 buffer[770] = 340;
 buffer[771] = 340;
 buffer[772] = 339;
 buffer[773] = 339;
 buffer[774] = 338;
 buffer[775] = 338;
 buffer[776] = 337;
 buffer[777] = 337;
 buffer[778] = 336;
 buffer[779] = 336;
 buffer[780] = 336;
 buffer[781] = 335;
 buffer[782] = 335;
 buffer[783] = 334;
 buffer[784] = 334;
 buffer[785] = 333;
 buffer[786] = 333;
 buffer[787] = 333;
 buffer[788] = 332;
 buffer[789] = 332;
 buffer[790] = 331;
 buffer[791] = 331;
 buffer[792] = 330;
 buffer[793] = 330;
 buffer[794] = 330;
 buffer[795] = 329;
 buffer[796] = 329;
 buffer[797] = 328;
 buffer[798] = 328;
 buffer[799] = 328;
 buffer[800] = 327;
 buffer[801] = 327;
 buffer[802] = 326;
 buffer[803] = 326;
 buffer[804] = 326;
 buffer[805] = 325;
 buffer[806] = 325;
 buffer[807] = 324;
 buffer[808] = 324;
 buffer[809] = 324;
 buffer[810] = 323;
 buffer[811] = 323;
 buffer[812] = 322;
 buffer[813] = 322;
 buffer[814] = 322;
 buffer[815] = 321;
 buffer[816] = 321;
 buffer[817] = 320;
 buffer[818] = 320;
 buffer[819] = 320;
 buffer[820] = 319;
 buffer[821] = 319;
 buffer[822] = 318;
 buffer[823] = 318;
 buffer[824] = 318;
 buffer[825] = 317;
 buffer[826] = 317;
 buffer[827] = 316;
 buffer[828] = 316;
 buffer[829] = 316;
 buffer[830] = 315;
 buffer[831] = 315;
 buffer[832] = 315;
 buffer[833] = 314;
 buffer[834] = 314;
 buffer[835] = 313;
 buffer[836] = 313;
 buffer[837] = 313;
 buffer[838] = 312;
 buffer[839] = 312;
 buffer[840] = 312;
 buffer[841] = 311;
 buffer[842] = 311;
 buffer[843] = 310;
 buffer[844] = 310;
 buffer[845] = 310;
 buffer[846] = 309;
 buffer[847] = 309;
 buffer[848] = 309;
 buffer[849] = 308;
 buffer[850] = 308;
 buffer[851] = 308;
 buffer[852] = 307;
 buffer[853] = 307;
 buffer[854] = 306;
 buffer[855] = 306;
 buffer[856] = 306;
 buffer[857] = 305;
 buffer[858] = 305;
 buffer[859] = 305;
 buffer[860] = 304;
 buffer[861] = 304;
 buffer[862] = 304;
 buffer[863] = 303;
 buffer[864] = 303;
 buffer[865] = 303;
 buffer[866] = 302;
 buffer[867] = 302;
 buffer[868] = 302;
 buffer[869] = 301;
 buffer[870] = 301;
 buffer[871] = 300;
 buffer[872] = 300;
 buffer[873] = 300;
 buffer[874] = 299;
 buffer[875] = 299;
 buffer[876] = 299;
 buffer[877] = 298;
 buffer[878] = 298;
 buffer[879] = 298;
 buffer[880] = 297;
 buffer[881] = 297;
 buffer[882] = 297;
 buffer[883] = 296;
 buffer[884] = 296;
 buffer[885] = 296;
 buffer[886] = 295;
 buffer[887] = 295;
 buffer[888] = 295;
 buffer[889] = 294;
 buffer[890] = 294;
 buffer[891] = 294;
 buffer[892] = 293;
 buffer[893] = 293;
 buffer[894] = 293;
 buffer[895] = 292;
 buffer[896] = 292;
 buffer[897] = 292;
 buffer[898] = 291;
 buffer[899] = 291;
 buffer[900] = 291;
 buffer[901] = 290;
 buffer[902] = 290;
 buffer[903] = 290;
 buffer[904] = 289;
 buffer[905] = 289;
 buffer[906] = 289;
 buffer[907] = 289;
 buffer[908] = 288;
 buffer[909] = 288;
 buffer[910] = 288;
 buffer[911] = 287;
 buffer[912] = 287;
 buffer[913] = 287;
 buffer[914] = 286;
 buffer[915] = 286;
 buffer[916] = 286;
 buffer[917] = 285;
 buffer[918] = 285;
 buffer[919] = 285;
 buffer[920] = 284;
 buffer[921] = 284;
 buffer[922] = 284;
 buffer[923] = 284;
 buffer[924] = 283;
 buffer[925] = 283;
 buffer[926] = 283;
 buffer[927] = 282;
 buffer[928] = 282;
 buffer[929] = 282;
 buffer[930] = 281;
 buffer[931] = 281;
 buffer[932] = 281;
 buffer[933] = 280;
 buffer[934] = 280;
 buffer[935] = 280;
 buffer[936] = 280;
 buffer[937] = 279;
 buffer[938] = 279;
 buffer[939] = 279;
 buffer[940] = 278;
 buffer[941] = 278;
 buffer[942] = 278;
 buffer[943] = 277;
 buffer[944] = 277;
 buffer[945] = 277;
 buffer[946] = 277;
 buffer[947] = 276;
 buffer[948] = 276;
 buffer[949] = 276;
 buffer[950] = 275;
 buffer[951] = 275;
 buffer[952] = 275;
 buffer[953] = 275;
 buffer[954] = 274;
 buffer[955] = 274;
 buffer[956] = 274;
 buffer[957] = 273;
 buffer[958] = 273;
 buffer[959] = 273;
 buffer[960] = 273;
 buffer[961] = 272;
 buffer[962] = 272;
 buffer[963] = 272;
 buffer[964] = 271;
 buffer[965] = 271;
 buffer[966] = 271;
 buffer[967] = 271;
 buffer[968] = 270;
 buffer[969] = 270;
 buffer[970] = 270;
 buffer[971] = 269;
 buffer[972] = 269;
 buffer[973] = 269;
 buffer[974] = 269;
 buffer[975] = 268;
 buffer[976] = 268;
 buffer[977] = 268;
 buffer[978] = 268;
 buffer[979] = 267;
 buffer[980] = 267;
 buffer[981] = 267;
 buffer[982] = 266;
 buffer[983] = 266;
 buffer[984] = 266;
 buffer[985] = 266;
 buffer[986] = 265;
 buffer[987] = 265;
 buffer[988] = 265;
 buffer[989] = 265;
 buffer[990] = 264;
 buffer[991] = 264;
 buffer[992] = 264;
 buffer[993] = 263;
 buffer[994] = 263;
 buffer[995] = 263;
 buffer[996] = 263;
 buffer[997] = 262;
 buffer[998] = 262;
 buffer[999] = 262;
 buffer[1000] = 262;
 buffer[1001] = 261;
 buffer[1002] = 261;
 buffer[1003] = 261;
 buffer[1004] = 261;
 buffer[1005] = 260;
 buffer[1006] = 260;
 buffer[1007] = 260;
 buffer[1008] = 260;
 buffer[1009] = 259;
 buffer[1010] = 259;
 buffer[1011] = 259;
 buffer[1012] = 259;
 buffer[1013] = 258;
 buffer[1014] = 258;
 buffer[1015] = 258;
 buffer[1016] = 258;
 buffer[1017] = 257;
 buffer[1018] = 257;
 buffer[1019] = 257;
 buffer[1020] = 257;
 buffer[1021] = 256;
 buffer[1022] = 256;
 buffer[1023] = 256;
 buffer[1024] = 256;
 buffer[1025] = 255;
 buffer[1026] = 255;
 buffer[1027] = 255;
 buffer[1028] = 255;
 buffer[1029] = 254;
 buffer[1030] = 254;
 buffer[1031] = 254;
 buffer[1032] = 254;
 buffer[1033] = 253;
 buffer[1034] = 253;
 buffer[1035] = 253;
 buffer[1036] = 253;
 buffer[1037] = 252;
 buffer[1038] = 252;
 buffer[1039] = 252;
 buffer[1040] = 252;
 buffer[1041] = 251;
 buffer[1042] = 251;
 buffer[1043] = 251;
 buffer[1044] = 251;
 buffer[1045] = 250;
 buffer[1046] = 250;
 buffer[1047] = 250;
 buffer[1048] = 250;
 buffer[1049] = 249;
 buffer[1050] = 249;
 buffer[1051] = 249;
 buffer[1052] = 249;
 buffer[1053] = 248;
 buffer[1054] = 248;
 buffer[1055] = 248;
 buffer[1056] = 248;
 buffer[1057] = 248;
 buffer[1058] = 247;
 buffer[1059] = 247;
 buffer[1060] = 247;
 buffer[1061] = 247;
 buffer[1062] = 246;
 buffer[1063] = 246;
 buffer[1064] = 246;
 buffer[1065] = 246;
 buffer[1066] = 245;
 buffer[1067] = 245;
 buffer[1068] = 245;
 buffer[1069] = 245;
 buffer[1070] = 244;
 buffer[1071] = 244;
 buffer[1072] = 244;
 buffer[1073] = 244;
 buffer[1074] = 244;
 buffer[1075] = 243;
 buffer[1076] = 243;
 buffer[1077] = 243;
 buffer[1078] = 243;
 buffer[1079] = 242;
 buffer[1080] = 242;
 buffer[1081] = 242;
 buffer[1082] = 242;
 buffer[1083] = 242;
 buffer[1084] = 241;
 buffer[1085] = 241;
 buffer[1086] = 241;
 buffer[1087] = 241;
 buffer[1088] = 240;
 buffer[1089] = 240;
 buffer[1090] = 240;
 buffer[1091] = 240;
 buffer[1092] = 240;
 buffer[1093] = 239;
 buffer[1094] = 239;
 buffer[1095] = 239;
 buffer[1096] = 239;
 buffer[1097] = 238;
 buffer[1098] = 238;
 buffer[1099] = 238;
 buffer[1100] = 238;
 buffer[1101] = 238;
 buffer[1102] = 237;
 buffer[1103] = 237;
 buffer[1104] = 237;
 buffer[1105] = 237;
 buffer[1106] = 237;
 buffer[1107] = 236;
 buffer[1108] = 236;
 buffer[1109] = 236;
 buffer[1110] = 236;
 buffer[1111] = 235;
 buffer[1112] = 235;
 buffer[1113] = 235;
 buffer[1114] = 235;
 buffer[1115] = 235;
 buffer[1116] = 234;
 buffer[1117] = 234;
 buffer[1118] = 234;
 buffer[1119] = 234;
 buffer[1120] = 234;
 buffer[1121] = 233;
 buffer[1122] = 233;
 buffer[1123] = 233;
 buffer[1124] = 233;
 buffer[1125] = 233;
 buffer[1126] = 232;
 buffer[1127] = 232;
 buffer[1128] = 232;
 buffer[1129] = 232;
 buffer[1130] = 231;
 buffer[1131] = 231;
 buffer[1132] = 231;
 buffer[1133] = 231;
 buffer[1134] = 231;
 buffer[1135] = 230;
 buffer[1136] = 230;
 buffer[1137] = 230;
 buffer[1138] = 230;
 buffer[1139] = 230;
 buffer[1140] = 229;
 buffer[1141] = 229;
 buffer[1142] = 229;
 buffer[1143] = 229;
 buffer[1144] = 229;
 buffer[1145] = 228;
 buffer[1146] = 228;
 buffer[1147] = 228;
 buffer[1148] = 228;
 buffer[1149] = 228;
 buffer[1150] = 227;
 buffer[1151] = 227;
 buffer[1152] = 227;
 buffer[1153] = 227;
 buffer[1154] = 227;
 buffer[1155] = 226;
 buffer[1156] = 226;
 buffer[1157] = 226;
 buffer[1158] = 226;
 buffer[1159] = 226;
 buffer[1160] = 225;
 buffer[1161] = 225;
 buffer[1162] = 225;
 buffer[1163] = 225;
 buffer[1164] = 225;
 buffer[1165] = 225;
 buffer[1166] = 224;
 buffer[1167] = 224;
 buffer[1168] = 224;
 buffer[1169] = 224;
 buffer[1170] = 224;
 buffer[1171] = 223;
 buffer[1172] = 223;
 buffer[1173] = 223;
 buffer[1174] = 223;
 buffer[1175] = 223;
 buffer[1176] = 222;
 buffer[1177] = 222;
 buffer[1178] = 222;
 buffer[1179] = 222;
 buffer[1180] = 222;
 buffer[1181] = 221;
 buffer[1182] = 221;
 buffer[1183] = 221;
 buffer[1184] = 221;
 buffer[1185] = 221;
 buffer[1186] = 221;
 buffer[1187] = 220;
 buffer[1188] = 220;
 buffer[1189] = 220;
 buffer[1190] = 220;
 buffer[1191] = 220;
 buffer[1192] = 219;
 buffer[1193] = 219;
 buffer[1194] = 219;
 buffer[1195] = 219;
 buffer[1196] = 219;
 buffer[1197] = 219;
 buffer[1198] = 218;
 buffer[1199] = 218;
 buffer[1200] = 218;
 buffer[1201] = 218;
 buffer[1202] = 218;
 buffer[1203] = 217;
 buffer[1204] = 217;
 buffer[1205] = 217;
 buffer[1206] = 217;
 buffer[1207] = 217;
 buffer[1208] = 217;
 buffer[1209] = 216;
 buffer[1210] = 216;
 buffer[1211] = 216;
 buffer[1212] = 216;
 buffer[1213] = 216;
 buffer[1214] = 215;
 buffer[1215] = 215;
 buffer[1216] = 215;
 buffer[1217] = 215;
 buffer[1218] = 215;
 buffer[1219] = 215;
 buffer[1220] = 214;
 buffer[1221] = 214;
 buffer[1222] = 214;
 buffer[1223] = 214;
 buffer[1224] = 214;
 buffer[1225] = 213;
 buffer[1226] = 213;
 buffer[1227] = 213;
 buffer[1228] = 213;
 buffer[1229] = 213;
 buffer[1230] = 213;
 buffer[1231] = 212;
 buffer[1232] = 212;
 buffer[1233] = 212;
 buffer[1234] = 212;
 buffer[1235] = 212;
 buffer[1236] = 212;
 buffer[1237] = 211;
 buffer[1238] = 211;
 buffer[1239] = 211;
 buffer[1240] = 211;
 buffer[1241] = 211;
 buffer[1242] = 211;
 buffer[1243] = 210;
 buffer[1244] = 210;
 buffer[1245] = 210;
 buffer[1246] = 210;
 buffer[1247] = 210;
 buffer[1248] = 210;
 buffer[1249] = 209;
 buffer[1250] = 209;
 buffer[1251] = 209;
 buffer[1252] = 209;
 buffer[1253] = 209;
 buffer[1254] = 209;
 buffer[1255] = 208;
 buffer[1256] = 208;
 buffer[1257] = 208;
 buffer[1258] = 208;
 buffer[1259] = 208;
 buffer[1260] = 208;
 buffer[1261] = 207;
 buffer[1262] = 207;
 buffer[1263] = 207;
 buffer[1264] = 207;
 buffer[1265] = 207;
 buffer[1266] = 207;
 buffer[1267] = 206;
 buffer[1268] = 206;
 buffer[1269] = 206;
 buffer[1270] = 206;
 buffer[1271] = 206;
 buffer[1272] = 206;
 buffer[1273] = 205;
 buffer[1274] = 205;
 buffer[1275] = 205;
 buffer[1276] = 205;
 buffer[1277] = 205;
 buffer[1278] = 205;
 buffer[1279] = 204;
 buffer[1280] = 204;
 buffer[1281] = 204;
 buffer[1282] = 204;
 buffer[1283] = 204;
 buffer[1284] = 204;
 buffer[1285] = 204;
 buffer[1286] = 203;
 buffer[1287] = 203;
 buffer[1288] = 203;
 buffer[1289] = 203;
 buffer[1290] = 203;
 buffer[1291] = 203;
 buffer[1292] = 202;
 buffer[1293] = 202;
 buffer[1294] = 202;
 buffer[1295] = 202;
 buffer[1296] = 202;
 buffer[1297] = 202;
 buffer[1298] = 201;
 buffer[1299] = 201;
 buffer[1300] = 201;
 buffer[1301] = 201;
 buffer[1302] = 201;
 buffer[1303] = 201;
 buffer[1304] = 201;
 buffer[1305] = 200;
 buffer[1306] = 200;
 buffer[1307] = 200;
 buffer[1308] = 200;
 buffer[1309] = 200;
 buffer[1310] = 200;
 buffer[1311] = 199;
 buffer[1312] = 199;
 buffer[1313] = 199;
 buffer[1314] = 199;
 buffer[1315] = 199;
 buffer[1316] = 199;
 buffer[1317] = 199;
 buffer[1318] = 198;
 buffer[1319] = 198;
 buffer[1320] = 198;
 buffer[1321] = 198;
 buffer[1322] = 198;
 buffer[1323] = 198;
 buffer[1324] = 197;
 buffer[1325] = 197;
 buffer[1326] = 197;
 buffer[1327] = 197;
 buffer[1328] = 197;
 buffer[1329] = 197;
 buffer[1330] = 197;
 buffer[1331] = 196;
 buffer[1332] = 196;
 buffer[1333] = 196;
 buffer[1334] = 196;
 buffer[1335] = 196;
 buffer[1336] = 196;
 buffer[1337] = 196;
 buffer[1338] = 195;
 buffer[1339] = 195;
 buffer[1340] = 195;
 buffer[1341] = 195;
 buffer[1342] = 195;
 buffer[1343] = 195;
 buffer[1344] = 195;
 buffer[1345] = 194;
 buffer[1346] = 194;
 buffer[1347] = 194;
 buffer[1348] = 194;
 buffer[1349] = 194;
 buffer[1350] = 194;
 buffer[1351] = 194;
 buffer[1352] = 193;
 buffer[1353] = 193;
 buffer[1354] = 193;
 buffer[1355] = 193;
 buffer[1356] = 193;
 buffer[1357] = 193;
 buffer[1358] = 193;
 buffer[1359] = 192;
 buffer[1360] = 192;
 buffer[1361] = 192;
 buffer[1362] = 192;
 buffer[1363] = 192;
 buffer[1364] = 192;
 buffer[1365] = 192;
 buffer[1366] = 191;
 buffer[1367] = 191;
 buffer[1368] = 191;
 buffer[1369] = 191;
 buffer[1370] = 191;
 buffer[1371] = 191;
 buffer[1372] = 191;
 buffer[1373] = 190;
 buffer[1374] = 190;
 buffer[1375] = 190;
 buffer[1376] = 190;
 buffer[1377] = 190;
 buffer[1378] = 190;
 buffer[1379] = 190;
 buffer[1380] = 189;
 buffer[1381] = 189;
 buffer[1382] = 189;
 buffer[1383] = 189;
 buffer[1384] = 189;
 buffer[1385] = 189;
 buffer[1386] = 189;
 buffer[1387] = 189;
 buffer[1388] = 188;
 buffer[1389] = 188;
 buffer[1390] = 188;
 buffer[1391] = 188;
 buffer[1392] = 188;
 buffer[1393] = 188;
 buffer[1394] = 188;
 buffer[1395] = 187;
 buffer[1396] = 187;
 buffer[1397] = 187;
 buffer[1398] = 187;
 buffer[1399] = 187;
 buffer[1400] = 187;
 buffer[1401] = 187;
 buffer[1402] = 186;
 buffer[1403] = 186;
 buffer[1404] = 186;
 buffer[1405] = 186;
 buffer[1406] = 186;
 buffer[1407] = 186;
 buffer[1408] = 186;
 buffer[1409] = 186;
 buffer[1410] = 185;
 buffer[1411] = 185;
 buffer[1412] = 185;
 buffer[1413] = 185;
 buffer[1414] = 185;
 buffer[1415] = 185;
 buffer[1416] = 185;
 buffer[1417] = 184;
 buffer[1418] = 184;
 buffer[1419] = 184;
 buffer[1420] = 184;
 buffer[1421] = 184;
 buffer[1422] = 184;
 buffer[1423] = 184;
 buffer[1424] = 184;
 buffer[1425] = 183;
 buffer[1426] = 183;
 buffer[1427] = 183;
 buffer[1428] = 183;
 buffer[1429] = 183;
 buffer[1430] = 183;
 buffer[1431] = 183;
 buffer[1432] = 183;
 buffer[1433] = 182;
 buffer[1434] = 182;
 buffer[1435] = 182;
 buffer[1436] = 182;
 buffer[1437] = 182;
 buffer[1438] = 182;
 buffer[1439] = 182;
 buffer[1440] = 182;
 buffer[1441] = 181;
 buffer[1442] = 181;
 buffer[1443] = 181;
 buffer[1444] = 181;
 buffer[1445] = 181;
 buffer[1446] = 181;
 buffer[1447] = 181;
 buffer[1448] = 181;
 buffer[1449] = 180;
 buffer[1450] = 180;
 buffer[1451] = 180;
 buffer[1452] = 180;
 buffer[1453] = 180;
 buffer[1454] = 180;
 buffer[1455] = 180;
 buffer[1456] = 180;
 buffer[1457] = 179;
 buffer[1458] = 179;
 buffer[1459] = 179;
 buffer[1460] = 179;
 buffer[1461] = 179;
 buffer[1462] = 179;
 buffer[1463] = 179;
 buffer[1464] = 179;
 buffer[1465] = 178;
 buffer[1466] = 178;
 buffer[1467] = 178;
 buffer[1468] = 178;
 buffer[1469] = 178;
 buffer[1470] = 178;
 buffer[1471] = 178;
 buffer[1472] = 178;
 buffer[1473] = 177;
 buffer[1474] = 177;
 buffer[1475] = 177;
 buffer[1476] = 177;
 buffer[1477] = 177;
 buffer[1478] = 177;
 buffer[1479] = 177;
 buffer[1480] = 177;
 buffer[1481] = 177;
 buffer[1482] = 176;
 buffer[1483] = 176;
 buffer[1484] = 176;
 buffer[1485] = 176;
 buffer[1486] = 176;
 buffer[1487] = 176;
 buffer[1488] = 176;
 buffer[1489] = 176;
 buffer[1490] = 175;
 buffer[1491] = 175;
 buffer[1492] = 175;
 buffer[1493] = 175;
 buffer[1494] = 175;
 buffer[1495] = 175;
 buffer[1496] = 175;
 buffer[1497] = 175;
 buffer[1498] = 174;
 buffer[1499] = 174;
 buffer[1500] = 174;
 buffer[1501] = 174;
 buffer[1502] = 174;
 buffer[1503] = 174;
 buffer[1504] = 174;
 buffer[1505] = 174;
 buffer[1506] = 174;
 buffer[1507] = 173;
 buffer[1508] = 173;
 buffer[1509] = 173;
 buffer[1510] = 173;
 buffer[1511] = 173;
 buffer[1512] = 173;
 buffer[1513] = 173;
 buffer[1514] = 173;
 buffer[1515] = 173;
 buffer[1516] = 172;
 buffer[1517] = 172;
 buffer[1518] = 172;
 buffer[1519] = 172;
 buffer[1520] = 172;
 buffer[1521] = 172;
 buffer[1522] = 172;
 buffer[1523] = 172;
 buffer[1524] = 172;
 buffer[1525] = 171;
 buffer[1526] = 171;
 buffer[1527] = 171;
 buffer[1528] = 171;
 buffer[1529] = 171;
 buffer[1530] = 171;
 buffer[1531] = 171;
 buffer[1532] = 171;
 buffer[1533] = 171;
 buffer[1534] = 170;
 buffer[1535] = 170;
 buffer[1536] = 170;
 buffer[1537] = 170;
 buffer[1538] = 170;
 buffer[1539] = 170;
 buffer[1540] = 170;
 buffer[1541] = 170;
 buffer[1542] = 170;
 buffer[1543] = 169;
 buffer[1544] = 169;
 buffer[1545] = 169;
 buffer[1546] = 169;
 buffer[1547] = 169;
 buffer[1548] = 169;
 buffer[1549] = 169;
 buffer[1550] = 169;
 buffer[1551] = 169;
 buffer[1552] = 168;
 buffer[1553] = 168;
 buffer[1554] = 168;
 buffer[1555] = 168;
 buffer[1556] = 168;
 buffer[1557] = 168;
 buffer[1558] = 168;
 buffer[1559] = 168;
 buffer[1560] = 168;
 buffer[1561] = 167;
 buffer[1562] = 167;
 buffer[1563] = 167;
 buffer[1564] = 167;
 buffer[1565] = 167;
 buffer[1566] = 167;
 buffer[1567] = 167;
 buffer[1568] = 167;
 buffer[1569] = 167;
 buffer[1570] = 166;
 buffer[1571] = 166;
 buffer[1572] = 166;
 buffer[1573] = 166;
 buffer[1574] = 166;
 buffer[1575] = 166;
 buffer[1576] = 166;
 buffer[1577] = 166;
 buffer[1578] = 166;
 buffer[1579] = 166;
 buffer[1580] = 165;
 buffer[1581] = 165;
 buffer[1582] = 165;
 buffer[1583] = 165;
 buffer[1584] = 165;
 buffer[1585] = 165;
 buffer[1586] = 165;
 buffer[1587] = 165;
 buffer[1588] = 165;
 buffer[1589] = 164;
 buffer[1590] = 164;
 buffer[1591] = 164;
 buffer[1592] = 164;
 buffer[1593] = 164;
 buffer[1594] = 164;
 buffer[1595] = 164;
 buffer[1596] = 164;
 buffer[1597] = 164;
 buffer[1598] = 164;
 buffer[1599] = 163;
 buffer[1600] = 163;
 buffer[1601] = 163;
 buffer[1602] = 163;
 buffer[1603] = 163;
 buffer[1604] = 163;
 buffer[1605] = 163;
 buffer[1606] = 163;
 buffer[1607] = 163;
 buffer[1608] = 163;
 buffer[1609] = 162;
 buffer[1610] = 162;
 buffer[1611] = 162;
 buffer[1612] = 162;
 buffer[1613] = 162;
 buffer[1614] = 162;
 buffer[1615] = 162;
 buffer[1616] = 162;
 buffer[1617] = 162;
 buffer[1618] = 162;
 buffer[1619] = 161;
 buffer[1620] = 161;
 buffer[1621] = 161;
 buffer[1622] = 161;
 buffer[1623] = 161;
 buffer[1624] = 161;
 buffer[1625] = 161;
 buffer[1626] = 161;
 buffer[1627] = 161;
 buffer[1628] = 161;
 buffer[1629] = 160;
 buffer[1630] = 160;
 buffer[1631] = 160;
 buffer[1632] = 160;
 buffer[1633] = 160;
 buffer[1634] = 160;
 buffer[1635] = 160;
 buffer[1636] = 160;
 buffer[1637] = 160;
 buffer[1638] = 160;
 buffer[1639] = 159;
 buffer[1640] = 159;
 buffer[1641] = 159;
 buffer[1642] = 159;
 buffer[1643] = 159;
 buffer[1644] = 159;
 buffer[1645] = 159;
 buffer[1646] = 159;
 buffer[1647] = 159;
 buffer[1648] = 159;
 buffer[1649] = 158;
 buffer[1650] = 158;
 buffer[1651] = 158;
 buffer[1652] = 158;
 buffer[1653] = 158;
 buffer[1654] = 158;
 buffer[1655] = 158;
 buffer[1656] = 158;
 buffer[1657] = 158;
 buffer[1658] = 158;
 buffer[1659] = 158;
 buffer[1660] = 157;
 buffer[1661] = 157;
 buffer[1662] = 157;
 buffer[1663] = 157;
 buffer[1664] = 157;
 buffer[1665] = 157;
 buffer[1666] = 157;
 buffer[1667] = 157;
 buffer[1668] = 157;
 buffer[1669] = 157;
 buffer[1670] = 156;
 buffer[1671] = 156;
 buffer[1672] = 156;
 buffer[1673] = 156;
 buffer[1674] = 156;
 buffer[1675] = 156;
 buffer[1676] = 156;
 buffer[1677] = 156;
 buffer[1678] = 156;
 buffer[1679] = 156;
 buffer[1680] = 156;
 buffer[1681] = 155;
 buffer[1682] = 155;
 buffer[1683] = 155;
 buffer[1684] = 155;
 buffer[1685] = 155;
 buffer[1686] = 155;
 buffer[1687] = 155;
 buffer[1688] = 155;
 buffer[1689] = 155;
 buffer[1690] = 155;
 buffer[1691] = 155;
 buffer[1692] = 154;
 buffer[1693] = 154;
 buffer[1694] = 154;
 buffer[1695] = 154;
 buffer[1696] = 154;
 buffer[1697] = 154;
 buffer[1698] = 154;
 buffer[1699] = 154;
 buffer[1700] = 154;
 buffer[1701] = 154;
 buffer[1702] = 154;
 buffer[1703] = 153;
 buffer[1704] = 153;
 buffer[1705] = 153;
 buffer[1706] = 153;
 buffer[1707] = 153;
 buffer[1708] = 153;
 buffer[1709] = 153;
 buffer[1710] = 153;
 buffer[1711] = 153;
 buffer[1712] = 153;
 buffer[1713] = 153;
 buffer[1714] = 152;
 buffer[1715] = 152;
 buffer[1716] = 152;
 buffer[1717] = 152;
 buffer[1718] = 152;
 buffer[1719] = 152;
 buffer[1720] = 152;
 buffer[1721] = 152;
 buffer[1722] = 152;
 buffer[1723] = 152;
 buffer[1724] = 152;
 buffer[1725] = 151;
 buffer[1726] = 151;
 buffer[1727] = 151;
 buffer[1728] = 151;
 buffer[1729] = 151;
 buffer[1730] = 151;
 buffer[1731] = 151;
 buffer[1732] = 151;
 buffer[1733] = 151;
 buffer[1734] = 151;
 buffer[1735] = 151;
 buffer[1736] = 151;
 buffer[1737] = 150;
 buffer[1738] = 150;
 buffer[1739] = 150;
 buffer[1740] = 150;
 buffer[1741] = 150;
 buffer[1742] = 150;
 buffer[1743] = 150;
 buffer[1744] = 150;
 buffer[1745] = 150;
 buffer[1746] = 150;
 buffer[1747] = 150;
 buffer[1748] = 149;
 buffer[1749] = 149;
 buffer[1750] = 149;
 buffer[1751] = 149;
 buffer[1752] = 149;
 buffer[1753] = 149;
 buffer[1754] = 149;
 buffer[1755] = 149;
 buffer[1756] = 149;
 buffer[1757] = 149;
 buffer[1758] = 149;
 buffer[1759] = 149;
 buffer[1760] = 148;
 buffer[1761] = 148;
 buffer[1762] = 148;
 buffer[1763] = 148;
 buffer[1764] = 148;
 buffer[1765] = 148;
 buffer[1766] = 148;
 buffer[1767] = 148;
 buffer[1768] = 148;
 buffer[1769] = 148;
 buffer[1770] = 148;
 buffer[1771] = 148;
 buffer[1772] = 147;
 buffer[1773] = 147;
 buffer[1774] = 147;
 buffer[1775] = 147;
 buffer[1776] = 147;
 buffer[1777] = 147;
 buffer[1778] = 147;
 buffer[1779] = 147;
 buffer[1780] = 147;
 buffer[1781] = 147;
 buffer[1782] = 147;
 buffer[1783] = 147;
 buffer[1784] = 146;
 buffer[1785] = 146;
 buffer[1786] = 146;
 buffer[1787] = 146;
 buffer[1788] = 146;
 buffer[1789] = 146;
 buffer[1790] = 146;
 buffer[1791] = 146;
 buffer[1792] = 146;
 buffer[1793] = 146;
 buffer[1794] = 146;
 buffer[1795] = 146;
 buffer[1796] = 145;
 buffer[1797] = 145;
 buffer[1798] = 145;
 buffer[1799] = 145;
 buffer[1800] = 145;
 buffer[1801] = 145;
 buffer[1802] = 145;
 buffer[1803] = 145;
 buffer[1804] = 145;
 buffer[1805] = 145;
 buffer[1806] = 145;
 buffer[1807] = 145;
 buffer[1808] = 144;
 buffer[1809] = 144;
 buffer[1810] = 144;
 buffer[1811] = 144;
 buffer[1812] = 144;
 buffer[1813] = 144;
 buffer[1814] = 144;
 buffer[1815] = 144;
 buffer[1816] = 144;
 buffer[1817] = 144;
 buffer[1818] = 144;
 buffer[1819] = 144;
 buffer[1820] = 144;
 buffer[1821] = 143;
 buffer[1822] = 143;
 buffer[1823] = 143;
 buffer[1824] = 143;
 buffer[1825] = 143;
 buffer[1826] = 143;
 buffer[1827] = 143;
 buffer[1828] = 143;
 buffer[1829] = 143;
 buffer[1830] = 143;
 buffer[1831] = 143;
 buffer[1832] = 143;
 buffer[1833] = 143;
 buffer[1834] = 142;
 buffer[1835] = 142;
 buffer[1836] = 142;
 buffer[1837] = 142;
 buffer[1838] = 142;
 buffer[1839] = 142;
 buffer[1840] = 142;
 buffer[1841] = 142;
 buffer[1842] = 142;
 buffer[1843] = 142;
 buffer[1844] = 142;
 buffer[1845] = 142;
 buffer[1846] = 142;
 buffer[1847] = 141;
 buffer[1848] = 141;
 buffer[1849] = 141;
 buffer[1850] = 141;
 buffer[1851] = 141;
 buffer[1852] = 141;
 buffer[1853] = 141;
 buffer[1854] = 141;
 buffer[1855] = 141;
 buffer[1856] = 141;
 buffer[1857] = 141;
 buffer[1858] = 141;
 buffer[1859] = 141;
 buffer[1860] = 140;
 buffer[1861] = 140;
 buffer[1862] = 140;
 buffer[1863] = 140;
 buffer[1864] = 140;
 buffer[1865] = 140;
 buffer[1866] = 140;
 buffer[1867] = 140;
 buffer[1868] = 140;
 buffer[1869] = 140;
 buffer[1870] = 140;
 buffer[1871] = 140;
 buffer[1872] = 140;
 buffer[1873] = 139;
 buffer[1874] = 139;
 buffer[1875] = 139;
 buffer[1876] = 139;
 buffer[1877] = 139;
 buffer[1878] = 139;
 buffer[1879] = 139;
 buffer[1880] = 139;
 buffer[1881] = 139;
 buffer[1882] = 139;
 buffer[1883] = 139;
 buffer[1884] = 139;
 buffer[1885] = 139;
 buffer[1886] = 138;
 buffer[1887] = 138;
 buffer[1888] = 138;
 buffer[1889] = 138;
 buffer[1890] = 138;
 buffer[1891] = 138;
 buffer[1892] = 138;
 buffer[1893] = 138;
 buffer[1894] = 138;
 buffer[1895] = 138;
 buffer[1896] = 138;
 buffer[1897] = 138;
 buffer[1898] = 138;
 buffer[1899] = 138;
 buffer[1900] = 137;
 buffer[1901] = 137;
 buffer[1902] = 137;
 buffer[1903] = 137;
 buffer[1904] = 137;
 buffer[1905] = 137;
 buffer[1906] = 137;
 buffer[1907] = 137;
 buffer[1908] = 137;
 buffer[1909] = 137;
 buffer[1910] = 137;
 buffer[1911] = 137;
 buffer[1912] = 137;
 buffer[1913] = 137;
 buffer[1914] = 136;
 buffer[1915] = 136;
 buffer[1916] = 136;
 buffer[1917] = 136;
 buffer[1918] = 136;
 buffer[1919] = 136;
 buffer[1920] = 136;
 buffer[1921] = 136;
 buffer[1922] = 136;
 buffer[1923] = 136;
 buffer[1924] = 136;
 buffer[1925] = 136;
 buffer[1926] = 136;
 buffer[1927] = 136;
 buffer[1928] = 135;
 buffer[1929] = 135;
 buffer[1930] = 135;
 buffer[1931] = 135;
 buffer[1932] = 135;
 buffer[1933] = 135;
 buffer[1934] = 135;
 buffer[1935] = 135;
 buffer[1936] = 135;
 buffer[1937] = 135;
 buffer[1938] = 135;
 buffer[1939] = 135;
 buffer[1940] = 135;
 buffer[1941] = 135;
 buffer[1942] = 134;
 buffer[1943] = 134;
 buffer[1944] = 134;
 buffer[1945] = 134;
 buffer[1946] = 134;
 buffer[1947] = 134;
 buffer[1948] = 134;
 buffer[1949] = 134;
 buffer[1950] = 134;
 buffer[1951] = 134;
 buffer[1952] = 134;
 buffer[1953] = 134;
 buffer[1954] = 134;
 buffer[1955] = 134;
 buffer[1956] = 134;
 buffer[1957] = 133;
 buffer[1958] = 133;
 buffer[1959] = 133;
 buffer[1960] = 133;
 buffer[1961] = 133;
 buffer[1962] = 133;
 buffer[1963] = 133;
 buffer[1964] = 133;
 buffer[1965] = 133;
 buffer[1966] = 133;
 buffer[1967] = 133;
 buffer[1968] = 133;
 buffer[1969] = 133;
 buffer[1970] = 133;
 buffer[1971] = 133;
 buffer[1972] = 132;
 buffer[1973] = 132;
 buffer[1974] = 132;
 buffer[1975] = 132;
 buffer[1976] = 132;
 buffer[1977] = 132;
 buffer[1978] = 132;
 buffer[1979] = 132;
 buffer[1980] = 132;
 buffer[1981] = 132;
 buffer[1982] = 132;
 buffer[1983] = 132;
 buffer[1984] = 132;
 buffer[1985] = 132;
 buffer[1986] = 131;
 buffer[1987] = 131;
 buffer[1988] = 131;
 buffer[1989] = 131;
 buffer[1990] = 131;
 buffer[1991] = 131;
 buffer[1992] = 131;
 buffer[1993] = 131;
 buffer[1994] = 131;
 buffer[1995] = 131;
 buffer[1996] = 131;
 buffer[1997] = 131;
 buffer[1998] = 131;
 buffer[1999] = 131;
 buffer[2000] = 131;
 buffer[2001] = 131;
 buffer[2002] = 130;
 buffer[2003] = 130;
 buffer[2004] = 130;
 buffer[2005] = 130;
 buffer[2006] = 130;
 buffer[2007] = 130;
 buffer[2008] = 130;
 buffer[2009] = 130;
 buffer[2010] = 130;
 buffer[2011] = 130;
 buffer[2012] = 130;
 buffer[2013] = 130;
 buffer[2014] = 130;
 buffer[2015] = 130;
 buffer[2016] = 130;
 buffer[2017] = 129;
 buffer[2018] = 129;
 buffer[2019] = 129;
 buffer[2020] = 129;
 buffer[2021] = 129;
 buffer[2022] = 129;
 buffer[2023] = 129;
 buffer[2024] = 129;
 buffer[2025] = 129;
 buffer[2026] = 129;
 buffer[2027] = 129;
 buffer[2028] = 129;
 buffer[2029] = 129;
 buffer[2030] = 129;
 buffer[2031] = 129;
 buffer[2032] = 129;
 buffer[2033] = 128;
 buffer[2034] = 128;
 buffer[2035] = 128;
 buffer[2036] = 128;
 buffer[2037] = 128;
 buffer[2038] = 128;
 buffer[2039] = 128;
 buffer[2040] = 128;
 buffer[2041] = 128;
 buffer[2042] = 128;
 buffer[2043] = 128;
 buffer[2044] = 128;
 buffer[2045] = 128;
 buffer[2046] = 128;
 buffer[2047] = 128;
end

endmodule

module M_frame_display (
in_pix_x,
in_pix_y,
in_pix_active,
in_pix_vblank,
in_vga_hs,
in_vga_vs,
out_pix_r,
out_pix_g,
out_pix_b,
in_run,
out_done,
reset,
out_clock,
clock
);
input  [10:0] in_pix_x;
input  [10:0] in_pix_y;
input  [0:0] in_pix_active;
input  [0:0] in_pix_vblank;
input  [0:0] in_vga_hs;
input  [0:0] in_vga_vs;
output  [7:0] out_pix_r;
output  [7:0] out_pix_g;
output  [7:0] out_pix_b;
input in_run;
output out_done;
input reset;
output out_clock;
input clock;
assign out_clock = clock;
wire signed [23:0] _w_mem_cos_rdata0;
wire signed [23:0] _w_mem_cos_rdata1;
wire signed [23:0] _w_mem_sin_rdata0;
wire signed [23:0] _w_mem_sin_rdata1;
wire  [17:0] _w_mem_invA_rdata0;
wire  [17:0] _w_mem_invA_rdata1;
wire  [17:0] _w_mem_invB_rdata;
wire signed [23:0] _c___stage___block_6_view_z;
assign _c___stage___block_6_view_z = 384;
wire  [0:0] _c___stage___block_6_inside;
assign _c___stage___block_6_inside = 0;
wire  [7:0] _c___stage___block_6_dist;
assign _c___stage___block_6_dist = 239;
wire  [7:0] _c___stage___block_6_clr;
assign _c___stage___block_6_clr = 0;
reg  [0:0] _t_cos_wenable0;
reg signed [23:0] _t_cos_wdata0;
reg  [0:0] _t_cos_wenable1;
reg signed [23:0] _t_cos_wdata1;
reg  [0:0] _t_sin_wenable0;
reg signed [23:0] _t_sin_wdata0;
reg  [0:0] _t_sin_wenable1;
reg signed [23:0] _t_sin_wdata1;
reg  [0:0] _t_invA_wenable0;
reg  [17:0] _t_invA_wdata0;
reg  [0:0] _t_invA_wenable1;
reg  [17:0] _t_invA_wdata1;
reg  [0:0] _t_invB_wenable;
reg  [17:0] _t_invB_wdata;
reg  [13:0] _t___stage___block_6_vxsz;
reg signed [23:0] _t___stage___block_6_view_x;
reg signed [23:0] _t___stage___block_6_view_y;
reg signed [23:0] _t___stage___block_7_cs0;
reg signed [23:0] _t___stage___block_7_ss0;
reg signed [23:0] _t___stage___block_7_cs1;
reg signed [23:0] _t___stage___block_7_ss1;
reg signed [23:0] _t___stage___block_7_rot_x;
reg signed [23:0] _t___stage___block_7_rot_y;
reg signed [23:0] _t___block_11_ycs;
reg signed [23:0] _t___block_11_yss;
reg signed [23:0] _t___stage___block_17_xcs;
reg signed [23:0] _t___block_19_xss;
reg signed [23:0] _t___block_21_zcs;
reg signed [23:0] _t___block_23_zss;
reg signed [23:0] _t___block_25_r_x_delta;
reg signed [23:0] _t___block_25_r_z_delta;
reg signed [15:0] _t___stage___block_26_rd_x;
reg signed [15:0] _t___stage___block_26_rd_y;
reg signed [15:0] _t___stage___block_26_rd_z;
reg signed [1:0] _t___stage___block_26_s_x;
reg signed [1:0] _t___stage___block_26_s_y;
reg signed [1:0] _t___stage___block_26_s_z;
reg signed [23:0] _t___stage___block_26_p_x;
reg signed [23:0] _t___stage___block_26_p_y;
reg signed [23:0] _t___stage___block_26_p_z;
reg signed [11:0] _t___stage___block_26_v_x;
reg signed [11:0] _t___stage___block_26_v_y;
reg signed [11:0] _t___stage___block_26_v_z;
reg  [13:0] _t___stage___block_26_brd_x;
reg  [13:0] _t___stage___block_26_brd_y;
reg  [13:0] _t___stage___block_26_brd_z;
reg  [17:0] _t___stage___block_28_inv_x;
reg  [17:0] _t___stage___block_28_inv_y;
reg  [17:0] _t___stage___block_28_inv_z;
reg  [31:0] _t___stage___block_28_tm_x_;
reg  [31:0] _t___stage___block_28_tm_y_;
reg  [31:0] _t___stage___block_28_tm_z_;
reg  [19:0] _t___block_34_tm_x;
reg  [19:0] _t___block_34_tm_y;
reg  [19:0] _t___block_34_tm_z;
reg  [31:0] _t___block_34_dt_x_;
reg  [31:0] _t___block_34_dt_y_;
reg  [31:0] _t___block_34_dt_z_;
reg  [19:0] _t___block_40_dt_x;
reg  [19:0] _t___block_40_dt_y;
reg  [19:0] _t___block_40_dt_z;
reg  [5:0] _t___stage___block_41_tex;
reg  [5:0] _t___stage___block_41_vnum0;
reg  [5:0] _t___stage___block_41_vnum1;
reg  [5:0] _t___stage___block_41_vnum2;
reg signed [20:0] _t___block_46_cmp_yx;
reg signed [20:0] _t___block_46_cmp_zx;
reg signed [20:0] _t___block_46_cmp_zy;
reg  [0:0] _t___block_46_x_sel;
reg  [0:0] _t___block_46_y_sel;
reg  [0:0] _t___block_46_z_sel;
reg  [5:0] _t___stage___block_62_tex;
reg  [5:0] _t___stage___block_62_vnum0;
reg  [5:0] _t___stage___block_62_vnum1;
reg  [5:0] _t___stage___block_62_vnum2;
reg signed [20:0] _t___block_67_cmp_yx;
reg signed [20:0] _t___block_67_cmp_zx;
reg signed [20:0] _t___block_67_cmp_zy;
reg  [0:0] _t___block_67_x_sel;
reg  [0:0] _t___block_67_y_sel;
reg  [0:0] _t___block_67_z_sel;
reg  [5:0] _t___stage___block_83_tex;
reg  [5:0] _t___stage___block_83_vnum0;
reg  [5:0] _t___stage___block_83_vnum1;
reg  [5:0] _t___stage___block_83_vnum2;
reg signed [20:0] _t___block_88_cmp_yx;
reg signed [20:0] _t___block_88_cmp_zx;
reg signed [20:0] _t___block_88_cmp_zy;
reg  [0:0] _t___block_88_x_sel;
reg  [0:0] _t___block_88_y_sel;
reg  [0:0] _t___block_88_z_sel;
reg  [5:0] _t___stage___block_104_tex;
reg  [5:0] _t___stage___block_104_vnum0;
reg  [5:0] _t___stage___block_104_vnum1;
reg  [5:0] _t___stage___block_104_vnum2;
reg signed [20:0] _t___block_109_cmp_yx;
reg signed [20:0] _t___block_109_cmp_zx;
reg signed [20:0] _t___block_109_cmp_zy;
reg  [0:0] _t___block_109_x_sel;
reg  [0:0] _t___block_109_y_sel;
reg  [0:0] _t___block_109_z_sel;
reg  [5:0] _t___stage___block_125_tex;
reg  [5:0] _t___stage___block_125_vnum0;
reg  [5:0] _t___stage___block_125_vnum1;
reg  [5:0] _t___stage___block_125_vnum2;
reg signed [20:0] _t___block_130_cmp_yx;
reg signed [20:0] _t___block_130_cmp_zx;
reg signed [20:0] _t___block_130_cmp_zy;
reg  [0:0] _t___block_130_x_sel;
reg  [0:0] _t___block_130_y_sel;
reg  [0:0] _t___block_130_z_sel;
reg  [5:0] _t___stage___block_146_tex;
reg  [5:0] _t___stage___block_146_vnum0;
reg  [5:0] _t___stage___block_146_vnum1;
reg  [5:0] _t___stage___block_146_vnum2;
reg signed [20:0] _t___block_151_cmp_yx;
reg signed [20:0] _t___block_151_cmp_zx;
reg signed [20:0] _t___block_151_cmp_zy;
reg  [0:0] _t___block_151_x_sel;
reg  [0:0] _t___block_151_y_sel;
reg  [0:0] _t___block_151_z_sel;
reg  [5:0] _t___stage___block_167_tex;
reg  [5:0] _t___stage___block_167_vnum0;
reg  [5:0] _t___stage___block_167_vnum1;
reg  [5:0] _t___stage___block_167_vnum2;
reg signed [20:0] _t___block_172_cmp_yx;
reg signed [20:0] _t___block_172_cmp_zx;
reg signed [20:0] _t___block_172_cmp_zy;
reg  [0:0] _t___block_172_x_sel;
reg  [0:0] _t___block_172_y_sel;
reg  [0:0] _t___block_172_z_sel;
reg  [5:0] _t___stage___block_188_tex;
reg  [5:0] _t___stage___block_188_vnum0;
reg  [5:0] _t___stage___block_188_vnum1;
reg  [5:0] _t___stage___block_188_vnum2;
reg signed [20:0] _t___block_193_cmp_yx;
reg signed [20:0] _t___block_193_cmp_zx;
reg signed [20:0] _t___block_193_cmp_zy;
reg  [0:0] _t___block_193_x_sel;
reg  [0:0] _t___block_193_y_sel;
reg  [0:0] _t___block_193_z_sel;
reg  [5:0] _t___stage___block_209_tex;
reg  [5:0] _t___stage___block_209_vnum0;
reg  [5:0] _t___stage___block_209_vnum1;
reg  [5:0] _t___stage___block_209_vnum2;
reg signed [20:0] _t___block_214_cmp_yx;
reg signed [20:0] _t___block_214_cmp_zx;
reg signed [20:0] _t___block_214_cmp_zy;
reg  [0:0] _t___block_214_x_sel;
reg  [0:0] _t___block_214_y_sel;
reg  [0:0] _t___block_214_z_sel;
reg  [5:0] _t___stage___block_230_tex;
reg  [5:0] _t___stage___block_230_vnum0;
reg  [5:0] _t___stage___block_230_vnum1;
reg  [5:0] _t___stage___block_230_vnum2;
reg signed [20:0] _t___block_235_cmp_yx;
reg signed [20:0] _t___block_235_cmp_zx;
reg signed [20:0] _t___block_235_cmp_zy;
reg  [0:0] _t___block_235_x_sel;
reg  [0:0] _t___block_235_y_sel;
reg  [0:0] _t___block_235_z_sel;
reg  [5:0] _t___stage___block_251_tex;
reg  [5:0] _t___stage___block_251_vnum0;
reg  [5:0] _t___stage___block_251_vnum1;
reg  [5:0] _t___stage___block_251_vnum2;
reg signed [20:0] _t___block_256_cmp_yx;
reg signed [20:0] _t___block_256_cmp_zx;
reg signed [20:0] _t___block_256_cmp_zy;
reg  [0:0] _t___block_256_x_sel;
reg  [0:0] _t___block_256_y_sel;
reg  [0:0] _t___block_256_z_sel;
reg  [5:0] _t___stage___block_272_tex;
reg  [5:0] _t___stage___block_272_vnum0;
reg  [5:0] _t___stage___block_272_vnum1;
reg  [5:0] _t___stage___block_272_vnum2;
reg signed [20:0] _t___block_277_cmp_yx;
reg signed [20:0] _t___block_277_cmp_zx;
reg signed [20:0] _t___block_277_cmp_zy;
reg  [0:0] _t___block_277_x_sel;
reg  [0:0] _t___block_277_y_sel;
reg  [0:0] _t___block_277_z_sel;
reg  [5:0] _t___stage___block_293_tex;
reg  [5:0] _t___stage___block_293_vnum0;
reg  [5:0] _t___stage___block_293_vnum1;
reg  [5:0] _t___stage___block_293_vnum2;
reg signed [20:0] _t___block_298_cmp_yx;
reg signed [20:0] _t___block_298_cmp_zx;
reg signed [20:0] _t___block_298_cmp_zy;
reg  [0:0] _t___block_298_x_sel;
reg  [0:0] _t___block_298_y_sel;
reg  [0:0] _t___block_298_z_sel;
reg  [5:0] _t___stage___block_314_tex;
reg  [5:0] _t___stage___block_314_vnum0;
reg  [5:0] _t___stage___block_314_vnum1;
reg  [5:0] _t___stage___block_314_vnum2;
reg signed [20:0] _t___block_319_cmp_yx;
reg signed [20:0] _t___block_319_cmp_zx;
reg signed [20:0] _t___block_319_cmp_zy;
reg  [0:0] _t___block_319_x_sel;
reg  [0:0] _t___block_319_y_sel;
reg  [0:0] _t___block_319_z_sel;
reg  [5:0] _t___stage___block_335_tex;
reg  [5:0] _t___stage___block_335_vnum0;
reg  [5:0] _t___stage___block_335_vnum1;
reg  [5:0] _t___stage___block_335_vnum2;
reg signed [20:0] _t___block_340_cmp_yx;
reg signed [20:0] _t___block_340_cmp_zx;
reg signed [20:0] _t___block_340_cmp_zy;
reg  [0:0] _t___block_340_x_sel;
reg  [0:0] _t___block_340_y_sel;
reg  [0:0] _t___block_340_z_sel;
reg  [5:0] _t___stage___block_356_tex;
reg  [5:0] _t___stage___block_356_vnum0;
reg  [5:0] _t___stage___block_356_vnum1;
reg  [5:0] _t___stage___block_356_vnum2;
reg signed [20:0] _t___block_361_cmp_yx;
reg signed [20:0] _t___block_361_cmp_zx;
reg signed [20:0] _t___block_361_cmp_zy;
reg  [0:0] _t___block_361_x_sel;
reg  [0:0] _t___block_361_y_sel;
reg  [0:0] _t___block_361_z_sel;
reg  [5:0] _t___stage___block_377_tex;
reg  [5:0] _t___stage___block_377_vnum0;
reg  [5:0] _t___stage___block_377_vnum1;
reg  [5:0] _t___stage___block_377_vnum2;
reg signed [20:0] _t___block_382_cmp_yx;
reg signed [20:0] _t___block_382_cmp_zx;
reg signed [20:0] _t___block_382_cmp_zy;
reg  [0:0] _t___block_382_x_sel;
reg  [0:0] _t___block_382_y_sel;
reg  [0:0] _t___block_382_z_sel;
reg  [5:0] _t___stage___block_398_tex;
reg  [5:0] _t___stage___block_398_vnum0;
reg  [5:0] _t___stage___block_398_vnum1;
reg  [5:0] _t___stage___block_398_vnum2;
reg signed [20:0] _t___block_403_cmp_yx;
reg signed [20:0] _t___block_403_cmp_zx;
reg signed [20:0] _t___block_403_cmp_zy;
reg  [0:0] _t___block_403_x_sel;
reg  [0:0] _t___block_403_y_sel;
reg  [0:0] _t___block_403_z_sel;
reg  [5:0] _t___stage___block_419_tex;
reg  [5:0] _t___stage___block_419_vnum0;
reg  [5:0] _t___stage___block_419_vnum1;
reg  [5:0] _t___stage___block_419_vnum2;
reg signed [20:0] _t___block_424_cmp_yx;
reg signed [20:0] _t___block_424_cmp_zx;
reg signed [20:0] _t___block_424_cmp_zy;
reg  [0:0] _t___block_424_x_sel;
reg  [0:0] _t___block_424_y_sel;
reg  [0:0] _t___block_424_z_sel;
reg  [5:0] _t___stage___block_440_tex;
reg  [5:0] _t___stage___block_440_vnum0;
reg  [5:0] _t___stage___block_440_vnum1;
reg  [5:0] _t___stage___block_440_vnum2;
reg signed [20:0] _t___block_445_cmp_yx;
reg signed [20:0] _t___block_445_cmp_zx;
reg signed [20:0] _t___block_445_cmp_zy;
reg  [0:0] _t___block_445_x_sel;
reg  [0:0] _t___block_445_y_sel;
reg  [0:0] _t___block_445_z_sel;
reg  [5:0] _t___stage___block_461_tex;
reg  [5:0] _t___stage___block_461_vnum0;
reg  [5:0] _t___stage___block_461_vnum1;
reg  [5:0] _t___stage___block_461_vnum2;
reg signed [20:0] _t___block_466_cmp_yx;
reg signed [20:0] _t___block_466_cmp_zx;
reg signed [20:0] _t___block_466_cmp_zy;
reg  [0:0] _t___block_466_x_sel;
reg  [0:0] _t___block_466_y_sel;
reg  [0:0] _t___block_466_z_sel;
reg  [5:0] _t___stage___block_482_tex;
reg  [5:0] _t___stage___block_482_vnum0;
reg  [5:0] _t___stage___block_482_vnum1;
reg  [5:0] _t___stage___block_482_vnum2;
reg signed [20:0] _t___block_487_cmp_yx;
reg signed [20:0] _t___block_487_cmp_zx;
reg signed [20:0] _t___block_487_cmp_zy;
reg  [0:0] _t___block_487_x_sel;
reg  [0:0] _t___block_487_y_sel;
reg  [0:0] _t___block_487_z_sel;
reg  [5:0] _t___stage___block_503_tex;
reg  [5:0] _t___stage___block_503_vnum0;
reg  [5:0] _t___stage___block_503_vnum1;
reg  [5:0] _t___stage___block_503_vnum2;
reg signed [20:0] _t___block_508_cmp_yx;
reg signed [20:0] _t___block_508_cmp_zx;
reg signed [20:0] _t___block_508_cmp_zy;
reg  [0:0] _t___block_508_x_sel;
reg  [0:0] _t___block_508_y_sel;
reg  [0:0] _t___block_508_z_sel;
reg  [5:0] _t___stage___block_524_tex;
reg  [5:0] _t___stage___block_524_vnum0;
reg  [5:0] _t___stage___block_524_vnum1;
reg  [5:0] _t___stage___block_524_vnum2;
reg signed [20:0] _t___block_529_cmp_yx;
reg signed [20:0] _t___block_529_cmp_zx;
reg signed [20:0] _t___block_529_cmp_zy;
reg  [0:0] _t___block_529_x_sel;
reg  [0:0] _t___block_529_y_sel;
reg  [0:0] _t___block_529_z_sel;
reg  [5:0] _t___stage___block_545_tex;
reg  [5:0] _t___stage___block_545_vnum0;
reg  [5:0] _t___stage___block_545_vnum1;
reg  [5:0] _t___stage___block_545_vnum2;
reg signed [20:0] _t___block_550_cmp_yx;
reg signed [20:0] _t___block_550_cmp_zx;
reg signed [20:0] _t___block_550_cmp_zy;
reg  [0:0] _t___block_550_x_sel;
reg  [0:0] _t___block_550_y_sel;
reg  [0:0] _t___block_550_z_sel;
reg  [5:0] _t___stage___block_566_tex;
reg  [5:0] _t___stage___block_566_vnum0;
reg  [5:0] _t___stage___block_566_vnum1;
reg  [5:0] _t___stage___block_566_vnum2;
reg signed [20:0] _t___block_571_cmp_yx;
reg signed [20:0] _t___block_571_cmp_zx;
reg signed [20:0] _t___block_571_cmp_zy;
reg  [0:0] _t___block_571_x_sel;
reg  [0:0] _t___block_571_y_sel;
reg  [0:0] _t___block_571_z_sel;
reg  [5:0] _t___stage___block_587_tex;
reg  [5:0] _t___stage___block_587_vnum0;
reg  [5:0] _t___stage___block_587_vnum1;
reg  [5:0] _t___stage___block_587_vnum2;
reg signed [20:0] _t___block_592_cmp_yx;
reg signed [20:0] _t___block_592_cmp_zx;
reg signed [20:0] _t___block_592_cmp_zy;
reg  [0:0] _t___block_592_x_sel;
reg  [0:0] _t___block_592_y_sel;
reg  [0:0] _t___block_592_z_sel;
reg  [5:0] _t___stage___block_608_tex;
reg  [5:0] _t___stage___block_608_vnum0;
reg  [5:0] _t___stage___block_608_vnum1;
reg  [5:0] _t___stage___block_608_vnum2;
reg signed [20:0] _t___block_613_cmp_yx;
reg signed [20:0] _t___block_613_cmp_zx;
reg signed [20:0] _t___block_613_cmp_zy;
reg  [0:0] _t___block_613_x_sel;
reg  [0:0] _t___block_613_y_sel;
reg  [0:0] _t___block_613_z_sel;
reg  [5:0] _t___stage___block_629_tex;
reg  [5:0] _t___stage___block_629_vnum0;
reg  [5:0] _t___stage___block_629_vnum1;
reg  [5:0] _t___stage___block_629_vnum2;
reg signed [20:0] _t___block_634_cmp_yx;
reg signed [20:0] _t___block_634_cmp_zx;
reg signed [20:0] _t___block_634_cmp_zy;
reg  [0:0] _t___block_634_x_sel;
reg  [0:0] _t___block_634_y_sel;
reg  [0:0] _t___block_634_z_sel;
reg  [5:0] _t___stage___block_650_tex;
reg  [5:0] _t___stage___block_650_vnum0;
reg  [5:0] _t___stage___block_650_vnum1;
reg  [5:0] _t___stage___block_650_vnum2;
reg signed [20:0] _t___block_655_cmp_yx;
reg signed [20:0] _t___block_655_cmp_zx;
reg signed [20:0] _t___block_655_cmp_zy;
reg  [0:0] _t___block_655_x_sel;
reg  [0:0] _t___block_655_y_sel;
reg  [0:0] _t___block_655_z_sel;
reg  [5:0] _t___stage___block_671_tex;
reg  [5:0] _t___stage___block_671_vnum0;
reg  [5:0] _t___stage___block_671_vnum1;
reg  [5:0] _t___stage___block_671_vnum2;
reg signed [20:0] _t___block_676_cmp_yx;
reg signed [20:0] _t___block_676_cmp_zx;
reg signed [20:0] _t___block_676_cmp_zy;
reg  [0:0] _t___block_676_x_sel;
reg  [0:0] _t___block_676_y_sel;
reg  [0:0] _t___block_676_z_sel;
reg  [5:0] _t___stage___block_692_tex;
reg  [5:0] _t___stage___block_692_vnum0;
reg  [5:0] _t___stage___block_692_vnum1;
reg  [5:0] _t___stage___block_692_vnum2;
reg signed [20:0] _t___block_697_cmp_yx;
reg signed [20:0] _t___block_697_cmp_zx;
reg signed [20:0] _t___block_697_cmp_zy;
reg  [0:0] _t___block_697_x_sel;
reg  [0:0] _t___block_697_y_sel;
reg  [0:0] _t___block_697_z_sel;
reg  [5:0] _t___stage___block_713_tex;
reg  [5:0] _t___stage___block_713_vnum0;
reg  [5:0] _t___stage___block_713_vnum1;
reg  [5:0] _t___stage___block_713_vnum2;
reg signed [20:0] _t___block_718_cmp_yx;
reg signed [20:0] _t___block_718_cmp_zx;
reg signed [20:0] _t___block_718_cmp_zy;
reg  [0:0] _t___block_718_x_sel;
reg  [0:0] _t___block_718_y_sel;
reg  [0:0] _t___block_718_z_sel;
reg  [5:0] _t___stage___block_734_tex;
reg  [5:0] _t___stage___block_734_vnum0;
reg  [5:0] _t___stage___block_734_vnum1;
reg  [5:0] _t___stage___block_734_vnum2;
reg signed [20:0] _t___block_739_cmp_yx;
reg signed [20:0] _t___block_739_cmp_zx;
reg signed [20:0] _t___block_739_cmp_zy;
reg  [0:0] _t___block_739_x_sel;
reg  [0:0] _t___block_739_y_sel;
reg  [0:0] _t___block_739_z_sel;
reg  [5:0] _t___stage___block_755_tex;
reg  [5:0] _t___stage___block_755_vnum0;
reg  [5:0] _t___stage___block_755_vnum1;
reg  [5:0] _t___stage___block_755_vnum2;
reg signed [20:0] _t___block_760_cmp_yx;
reg signed [20:0] _t___block_760_cmp_zx;
reg signed [20:0] _t___block_760_cmp_zy;
reg  [0:0] _t___block_760_x_sel;
reg  [0:0] _t___block_760_y_sel;
reg  [0:0] _t___block_760_z_sel;
reg  [5:0] _t___stage___block_776_tex;
reg  [5:0] _t___stage___block_776_vnum0;
reg  [5:0] _t___stage___block_776_vnum1;
reg  [5:0] _t___stage___block_776_vnum2;
reg signed [20:0] _t___block_781_cmp_yx;
reg signed [20:0] _t___block_781_cmp_zx;
reg signed [20:0] _t___block_781_cmp_zy;
reg  [0:0] _t___block_781_x_sel;
reg  [0:0] _t___block_781_y_sel;
reg  [0:0] _t___block_781_z_sel;
reg  [5:0] _t___stage___block_797_tex;
reg  [5:0] _t___stage___block_797_vnum0;
reg  [5:0] _t___stage___block_797_vnum1;
reg  [5:0] _t___stage___block_797_vnum2;
reg signed [20:0] _t___block_802_cmp_yx;
reg signed [20:0] _t___block_802_cmp_zx;
reg signed [20:0] _t___block_802_cmp_zy;
reg  [0:0] _t___block_802_x_sel;
reg  [0:0] _t___block_802_y_sel;
reg  [0:0] _t___block_802_z_sel;
reg  [5:0] _t___stage___block_818_tex;
reg  [5:0] _t___stage___block_818_vnum0;
reg  [5:0] _t___stage___block_818_vnum1;
reg  [5:0] _t___stage___block_818_vnum2;
reg signed [20:0] _t___block_823_cmp_yx;
reg signed [20:0] _t___block_823_cmp_zx;
reg signed [20:0] _t___block_823_cmp_zy;
reg  [0:0] _t___block_823_x_sel;
reg  [0:0] _t___block_823_y_sel;
reg  [0:0] _t___block_823_z_sel;
reg  [5:0] _t___stage___block_839_tex;
reg  [5:0] _t___stage___block_839_vnum0;
reg  [5:0] _t___stage___block_839_vnum1;
reg  [5:0] _t___stage___block_839_vnum2;
reg signed [20:0] _t___block_844_cmp_yx;
reg signed [20:0] _t___block_844_cmp_zx;
reg signed [20:0] _t___block_844_cmp_zy;
reg  [0:0] _t___block_844_x_sel;
reg  [0:0] _t___block_844_y_sel;
reg  [0:0] _t___block_844_z_sel;
reg  [5:0] _t___stage___block_860_tex;
reg  [5:0] _t___stage___block_860_vnum0;
reg  [5:0] _t___stage___block_860_vnum1;
reg  [5:0] _t___stage___block_860_vnum2;
reg signed [20:0] _t___block_865_cmp_yx;
reg signed [20:0] _t___block_865_cmp_zx;
reg signed [20:0] _t___block_865_cmp_zy;
reg  [0:0] _t___block_865_x_sel;
reg  [0:0] _t___block_865_y_sel;
reg  [0:0] _t___block_865_z_sel;
reg  [5:0] _t___stage___block_881_tex;
reg  [5:0] _t___stage___block_881_vnum0;
reg  [5:0] _t___stage___block_881_vnum1;
reg  [5:0] _t___stage___block_881_vnum2;
reg signed [20:0] _t___block_886_cmp_yx;
reg signed [20:0] _t___block_886_cmp_zx;
reg signed [20:0] _t___block_886_cmp_zy;
reg  [0:0] _t___block_886_x_sel;
reg  [0:0] _t___block_886_y_sel;
reg  [0:0] _t___block_886_z_sel;
reg  [5:0] _t___stage___block_902_tex;
reg  [5:0] _t___stage___block_902_vnum0;
reg  [5:0] _t___stage___block_902_vnum1;
reg  [5:0] _t___stage___block_902_vnum2;
reg signed [20:0] _t___block_907_cmp_yx;
reg signed [20:0] _t___block_907_cmp_zx;
reg signed [20:0] _t___block_907_cmp_zy;
reg  [0:0] _t___block_907_x_sel;
reg  [0:0] _t___block_907_y_sel;
reg  [0:0] _t___block_907_z_sel;
reg  [5:0] _t___stage___block_923_tex;
reg  [5:0] _t___stage___block_923_vnum0;
reg  [5:0] _t___stage___block_923_vnum1;
reg  [5:0] _t___stage___block_923_vnum2;
reg signed [20:0] _t___block_928_cmp_yx;
reg signed [20:0] _t___block_928_cmp_zx;
reg signed [20:0] _t___block_928_cmp_zy;
reg  [0:0] _t___block_928_x_sel;
reg  [0:0] _t___block_928_y_sel;
reg  [0:0] _t___block_928_z_sel;
reg  [5:0] _t___stage___block_944_tex;
reg  [5:0] _t___stage___block_944_vnum0;
reg  [5:0] _t___stage___block_944_vnum1;
reg  [5:0] _t___stage___block_944_vnum2;
reg signed [20:0] _t___block_949_cmp_yx;
reg signed [20:0] _t___block_949_cmp_zx;
reg signed [20:0] _t___block_949_cmp_zy;
reg  [0:0] _t___block_949_x_sel;
reg  [0:0] _t___block_949_y_sel;
reg  [0:0] _t___block_949_z_sel;
reg  [5:0] _t___stage___block_965_tex;
reg  [5:0] _t___stage___block_965_vnum0;
reg  [5:0] _t___stage___block_965_vnum1;
reg  [5:0] _t___stage___block_965_vnum2;
reg signed [20:0] _t___block_970_cmp_yx;
reg signed [20:0] _t___block_970_cmp_zx;
reg signed [20:0] _t___block_970_cmp_zy;
reg  [0:0] _t___block_970_x_sel;
reg  [0:0] _t___block_970_y_sel;
reg  [0:0] _t___block_970_z_sel;
reg  [5:0] _t___stage___block_986_tex;
reg  [5:0] _t___stage___block_986_vnum0;
reg  [5:0] _t___stage___block_986_vnum1;
reg  [5:0] _t___stage___block_986_vnum2;
reg signed [20:0] _t___block_991_cmp_yx;
reg signed [20:0] _t___block_991_cmp_zx;
reg signed [20:0] _t___block_991_cmp_zy;
reg  [0:0] _t___block_991_x_sel;
reg  [0:0] _t___block_991_y_sel;
reg  [0:0] _t___block_991_z_sel;
reg  [5:0] _t___stage___block_1007_tex;
reg  [5:0] _t___stage___block_1007_vnum0;
reg  [5:0] _t___stage___block_1007_vnum1;
reg  [5:0] _t___stage___block_1007_vnum2;
reg signed [20:0] _t___block_1012_cmp_yx;
reg signed [20:0] _t___block_1012_cmp_zx;
reg signed [20:0] _t___block_1012_cmp_zy;
reg  [0:0] _t___block_1012_x_sel;
reg  [0:0] _t___block_1012_y_sel;
reg  [0:0] _t___block_1012_z_sel;
reg  [5:0] _t___stage___block_1028_tex;
reg  [5:0] _t___stage___block_1028_vnum0;
reg  [5:0] _t___stage___block_1028_vnum1;
reg  [5:0] _t___stage___block_1028_vnum2;
reg signed [20:0] _t___block_1033_cmp_yx;
reg signed [20:0] _t___block_1033_cmp_zx;
reg signed [20:0] _t___block_1033_cmp_zy;
reg  [0:0] _t___block_1033_x_sel;
reg  [0:0] _t___block_1033_y_sel;
reg  [0:0] _t___block_1033_z_sel;
reg  [5:0] _t___stage___block_1049_tex;
reg  [5:0] _t___stage___block_1049_vnum0;
reg  [5:0] _t___stage___block_1049_vnum1;
reg  [5:0] _t___stage___block_1049_vnum2;
reg signed [20:0] _t___block_1054_cmp_yx;
reg signed [20:0] _t___block_1054_cmp_zx;
reg signed [20:0] _t___block_1054_cmp_zy;
reg  [0:0] _t___block_1054_x_sel;
reg  [0:0] _t___block_1054_y_sel;
reg  [0:0] _t___block_1054_z_sel;
reg  [5:0] _t___stage___block_1070_tex;
reg  [5:0] _t___stage___block_1070_vnum0;
reg  [5:0] _t___stage___block_1070_vnum1;
reg  [5:0] _t___stage___block_1070_vnum2;
reg signed [20:0] _t___block_1075_cmp_yx;
reg signed [20:0] _t___block_1075_cmp_zx;
reg signed [20:0] _t___block_1075_cmp_zy;
reg  [0:0] _t___block_1075_x_sel;
reg  [0:0] _t___block_1075_y_sel;
reg  [0:0] _t___block_1075_z_sel;
reg  [5:0] _t___stage___block_1091_tex;
reg  [5:0] _t___stage___block_1091_vnum0;
reg  [5:0] _t___stage___block_1091_vnum1;
reg  [5:0] _t___stage___block_1091_vnum2;
reg signed [20:0] _t___block_1096_cmp_yx;
reg signed [20:0] _t___block_1096_cmp_zx;
reg signed [20:0] _t___block_1096_cmp_zy;
reg  [0:0] _t___block_1096_x_sel;
reg  [0:0] _t___block_1096_y_sel;
reg  [0:0] _t___block_1096_z_sel;
reg  [5:0] _t___stage___block_1112_tex;
reg  [5:0] _t___stage___block_1112_vnum0;
reg  [5:0] _t___stage___block_1112_vnum1;
reg  [5:0] _t___stage___block_1112_vnum2;
reg signed [20:0] _t___block_1117_cmp_yx;
reg signed [20:0] _t___block_1117_cmp_zx;
reg signed [20:0] _t___block_1117_cmp_zy;
reg  [0:0] _t___block_1117_x_sel;
reg  [0:0] _t___block_1117_y_sel;
reg  [0:0] _t___block_1117_z_sel;
reg  [5:0] _t___stage___block_1133_tex;
reg  [5:0] _t___stage___block_1133_vnum0;
reg  [5:0] _t___stage___block_1133_vnum1;
reg  [5:0] _t___stage___block_1133_vnum2;
reg signed [20:0] _t___block_1138_cmp_yx;
reg signed [20:0] _t___block_1138_cmp_zx;
reg signed [20:0] _t___block_1138_cmp_zy;
reg  [0:0] _t___block_1138_x_sel;
reg  [0:0] _t___block_1138_y_sel;
reg  [0:0] _t___block_1138_z_sel;
reg  [5:0] _t___stage___block_1154_tex;
reg  [5:0] _t___stage___block_1154_vnum0;
reg  [5:0] _t___stage___block_1154_vnum1;
reg  [5:0] _t___stage___block_1154_vnum2;
reg signed [20:0] _t___block_1159_cmp_yx;
reg signed [20:0] _t___block_1159_cmp_zx;
reg signed [20:0] _t___block_1159_cmp_zy;
reg  [0:0] _t___block_1159_x_sel;
reg  [0:0] _t___block_1159_y_sel;
reg  [0:0] _t___block_1159_z_sel;
reg  [5:0] _t___stage___block_1175_tex;
reg  [5:0] _t___stage___block_1175_vnum0;
reg  [5:0] _t___stage___block_1175_vnum1;
reg  [5:0] _t___stage___block_1175_vnum2;
reg signed [20:0] _t___block_1180_cmp_yx;
reg signed [20:0] _t___block_1180_cmp_zx;
reg signed [20:0] _t___block_1180_cmp_zy;
reg  [0:0] _t___block_1180_x_sel;
reg  [0:0] _t___block_1180_y_sel;
reg  [0:0] _t___block_1180_z_sel;
reg  [5:0] _t___stage___block_1196_tex;
reg  [5:0] _t___stage___block_1196_vnum0;
reg  [5:0] _t___stage___block_1196_vnum1;
reg  [5:0] _t___stage___block_1196_vnum2;
reg signed [20:0] _t___block_1201_cmp_yx;
reg signed [20:0] _t___block_1201_cmp_zx;
reg signed [20:0] _t___block_1201_cmp_zy;
reg  [0:0] _t___block_1201_x_sel;
reg  [0:0] _t___block_1201_y_sel;
reg  [0:0] _t___block_1201_z_sel;
reg  [5:0] _t___stage___block_1217_tex;
reg  [5:0] _t___stage___block_1217_vnum0;
reg  [5:0] _t___stage___block_1217_vnum1;
reg  [5:0] _t___stage___block_1217_vnum2;
reg signed [20:0] _t___block_1222_cmp_yx;
reg signed [20:0] _t___block_1222_cmp_zx;
reg signed [20:0] _t___block_1222_cmp_zy;
reg  [0:0] _t___block_1222_x_sel;
reg  [0:0] _t___block_1222_y_sel;
reg  [0:0] _t___block_1222_z_sel;
reg  [5:0] _t___stage___block_1238_tex;
reg  [5:0] _t___stage___block_1238_vnum0;
reg  [5:0] _t___stage___block_1238_vnum1;
reg  [5:0] _t___stage___block_1238_vnum2;
reg signed [20:0] _t___block_1243_cmp_yx;
reg signed [20:0] _t___block_1243_cmp_zx;
reg signed [20:0] _t___block_1243_cmp_zy;
reg  [0:0] _t___block_1243_x_sel;
reg  [0:0] _t___block_1243_y_sel;
reg  [0:0] _t___block_1243_z_sel;
reg  [5:0] _t___stage___block_1259_tex;
reg  [5:0] _t___stage___block_1259_vnum0;
reg  [5:0] _t___stage___block_1259_vnum1;
reg  [5:0] _t___stage___block_1259_vnum2;
reg signed [20:0] _t___block_1264_cmp_yx;
reg signed [20:0] _t___block_1264_cmp_zx;
reg signed [20:0] _t___block_1264_cmp_zy;
reg  [0:0] _t___block_1264_x_sel;
reg  [0:0] _t___block_1264_y_sel;
reg  [0:0] _t___block_1264_z_sel;
reg  [5:0] _t___stage___block_1280_tex;
reg  [5:0] _t___stage___block_1280_vnum0;
reg  [5:0] _t___stage___block_1280_vnum1;
reg  [5:0] _t___stage___block_1280_vnum2;
reg signed [20:0] _t___block_1285_cmp_yx;
reg signed [20:0] _t___block_1285_cmp_zx;
reg signed [20:0] _t___block_1285_cmp_zy;
reg  [0:0] _t___block_1285_x_sel;
reg  [0:0] _t___block_1285_y_sel;
reg  [0:0] _t___block_1285_z_sel;
reg  [5:0] _t___stage___block_1301_tex;
reg  [5:0] _t___stage___block_1301_vnum0;
reg  [5:0] _t___stage___block_1301_vnum1;
reg  [5:0] _t___stage___block_1301_vnum2;
reg signed [20:0] _t___block_1306_cmp_yx;
reg signed [20:0] _t___block_1306_cmp_zx;
reg signed [20:0] _t___block_1306_cmp_zy;
reg  [0:0] _t___block_1306_x_sel;
reg  [0:0] _t___block_1306_y_sel;
reg  [0:0] _t___block_1306_z_sel;
reg  [5:0] _t___stage___block_1322_tex;
reg  [5:0] _t___stage___block_1322_vnum0;
reg  [5:0] _t___stage___block_1322_vnum1;
reg  [5:0] _t___stage___block_1322_vnum2;
reg signed [20:0] _t___block_1327_cmp_yx;
reg signed [20:0] _t___block_1327_cmp_zx;
reg signed [20:0] _t___block_1327_cmp_zy;
reg  [0:0] _t___block_1327_x_sel;
reg  [0:0] _t___block_1327_y_sel;
reg  [0:0] _t___block_1327_z_sel;
reg  [5:0] _t___stage___block_1343_tex;
reg  [5:0] _t___stage___block_1343_vnum0;
reg  [5:0] _t___stage___block_1343_vnum1;
reg  [5:0] _t___stage___block_1343_vnum2;
reg signed [20:0] _t___block_1348_cmp_yx;
reg signed [20:0] _t___block_1348_cmp_zx;
reg signed [20:0] _t___block_1348_cmp_zy;
reg  [0:0] _t___block_1348_x_sel;
reg  [0:0] _t___block_1348_y_sel;
reg  [0:0] _t___block_1348_z_sel;
reg  [5:0] _t___stage___block_1364_tex;
reg  [5:0] _t___stage___block_1364_vnum0;
reg  [5:0] _t___stage___block_1364_vnum1;
reg  [5:0] _t___stage___block_1364_vnum2;
reg signed [20:0] _t___block_1369_cmp_yx;
reg signed [20:0] _t___block_1369_cmp_zx;
reg signed [20:0] _t___block_1369_cmp_zy;
reg  [0:0] _t___block_1369_x_sel;
reg  [0:0] _t___block_1369_y_sel;
reg  [0:0] _t___block_1369_z_sel;
reg  [5:0] _t___stage___block_1385_tex;
reg  [5:0] _t___stage___block_1385_vnum0;
reg  [5:0] _t___stage___block_1385_vnum1;
reg  [5:0] _t___stage___block_1385_vnum2;
reg signed [20:0] _t___block_1390_cmp_yx;
reg signed [20:0] _t___block_1390_cmp_zx;
reg signed [20:0] _t___block_1390_cmp_zy;
reg  [0:0] _t___block_1390_x_sel;
reg  [0:0] _t___block_1390_y_sel;
reg  [0:0] _t___block_1390_z_sel;
reg  [5:0] _t___stage___block_1406_tex;
reg  [5:0] _t___stage___block_1406_vnum0;
reg  [5:0] _t___stage___block_1406_vnum1;
reg  [5:0] _t___stage___block_1406_vnum2;
reg signed [20:0] _t___block_1411_cmp_yx;
reg signed [20:0] _t___block_1411_cmp_zx;
reg signed [20:0] _t___block_1411_cmp_zy;
reg  [0:0] _t___block_1411_x_sel;
reg  [0:0] _t___block_1411_y_sel;
reg  [0:0] _t___block_1411_z_sel;
reg  [5:0] _t___stage___block_1427_tex;
reg  [5:0] _t___stage___block_1427_vnum0;
reg  [5:0] _t___stage___block_1427_vnum1;
reg  [5:0] _t___stage___block_1427_vnum2;
reg signed [20:0] _t___block_1432_cmp_yx;
reg signed [20:0] _t___block_1432_cmp_zx;
reg signed [20:0] _t___block_1432_cmp_zy;
reg  [0:0] _t___block_1432_x_sel;
reg  [0:0] _t___block_1432_y_sel;
reg  [0:0] _t___block_1432_z_sel;
reg  [5:0] _t___stage___block_1448_tex;
reg  [5:0] _t___stage___block_1448_vnum0;
reg  [5:0] _t___stage___block_1448_vnum1;
reg  [5:0] _t___stage___block_1448_vnum2;
reg signed [20:0] _t___block_1453_cmp_yx;
reg signed [20:0] _t___block_1453_cmp_zx;
reg signed [20:0] _t___block_1453_cmp_zy;
reg  [0:0] _t___block_1453_x_sel;
reg  [0:0] _t___block_1453_y_sel;
reg  [0:0] _t___block_1453_z_sel;
reg  [5:0] _t___stage___block_1469_tex;
reg  [5:0] _t___stage___block_1469_vnum0;
reg  [5:0] _t___stage___block_1469_vnum1;
reg  [5:0] _t___stage___block_1469_vnum2;
reg signed [20:0] _t___block_1474_cmp_yx;
reg signed [20:0] _t___block_1474_cmp_zx;
reg signed [20:0] _t___block_1474_cmp_zy;
reg  [0:0] _t___block_1474_x_sel;
reg  [0:0] _t___block_1474_y_sel;
reg  [0:0] _t___block_1474_z_sel;
reg  [5:0] _t___stage___block_1490_tex;
reg  [5:0] _t___stage___block_1490_vnum0;
reg  [5:0] _t___stage___block_1490_vnum1;
reg  [5:0] _t___stage___block_1490_vnum2;
reg signed [20:0] _t___block_1495_cmp_yx;
reg signed [20:0] _t___block_1495_cmp_zx;
reg signed [20:0] _t___block_1495_cmp_zy;
reg  [0:0] _t___block_1495_x_sel;
reg  [0:0] _t___block_1495_y_sel;
reg  [0:0] _t___block_1495_z_sel;
reg  [5:0] _t___stage___block_1511_tex;
reg  [5:0] _t___stage___block_1511_vnum0;
reg  [5:0] _t___stage___block_1511_vnum1;
reg  [5:0] _t___stage___block_1511_vnum2;
reg signed [20:0] _t___block_1516_cmp_yx;
reg signed [20:0] _t___block_1516_cmp_zx;
reg signed [20:0] _t___block_1516_cmp_zy;
reg  [0:0] _t___block_1516_x_sel;
reg  [0:0] _t___block_1516_y_sel;
reg  [0:0] _t___block_1516_z_sel;
reg  [5:0] _t___stage___block_1532_tex;
reg  [5:0] _t___stage___block_1532_vnum0;
reg  [5:0] _t___stage___block_1532_vnum1;
reg  [5:0] _t___stage___block_1532_vnum2;
reg signed [20:0] _t___block_1537_cmp_yx;
reg signed [20:0] _t___block_1537_cmp_zx;
reg signed [20:0] _t___block_1537_cmp_zy;
reg  [0:0] _t___block_1537_x_sel;
reg  [0:0] _t___block_1537_y_sel;
reg  [0:0] _t___block_1537_z_sel;
reg  [5:0] _t___stage___block_1553_tex;
reg  [5:0] _t___stage___block_1553_vnum0;
reg  [5:0] _t___stage___block_1553_vnum1;
reg  [5:0] _t___stage___block_1553_vnum2;
reg signed [20:0] _t___block_1558_cmp_yx;
reg signed [20:0] _t___block_1558_cmp_zx;
reg signed [20:0] _t___block_1558_cmp_zy;
reg  [0:0] _t___block_1558_x_sel;
reg  [0:0] _t___block_1558_y_sel;
reg  [0:0] _t___block_1558_z_sel;
reg  [5:0] _t___stage___block_1574_tex;
reg  [5:0] _t___stage___block_1574_vnum0;
reg  [5:0] _t___stage___block_1574_vnum1;
reg  [5:0] _t___stage___block_1574_vnum2;
reg signed [20:0] _t___block_1579_cmp_yx;
reg signed [20:0] _t___block_1579_cmp_zx;
reg signed [20:0] _t___block_1579_cmp_zy;
reg  [0:0] _t___block_1579_x_sel;
reg  [0:0] _t___block_1579_y_sel;
reg  [0:0] _t___block_1579_z_sel;
reg  [5:0] _t___stage___block_1595_tex;
reg  [5:0] _t___stage___block_1595_vnum0;
reg  [5:0] _t___stage___block_1595_vnum1;
reg  [5:0] _t___stage___block_1595_vnum2;
reg signed [20:0] _t___block_1600_cmp_yx;
reg signed [20:0] _t___block_1600_cmp_zx;
reg signed [20:0] _t___block_1600_cmp_zy;
reg  [0:0] _t___block_1600_x_sel;
reg  [0:0] _t___block_1600_y_sel;
reg  [0:0] _t___block_1600_z_sel;
reg  [5:0] _t___stage___block_1616_tex;
reg  [5:0] _t___stage___block_1616_vnum0;
reg  [5:0] _t___stage___block_1616_vnum1;
reg  [5:0] _t___stage___block_1616_vnum2;
reg signed [20:0] _t___block_1621_cmp_yx;
reg signed [20:0] _t___block_1621_cmp_zx;
reg signed [20:0] _t___block_1621_cmp_zy;
reg  [0:0] _t___block_1621_x_sel;
reg  [0:0] _t___block_1621_y_sel;
reg  [0:0] _t___block_1621_z_sel;
reg  [5:0] _t___stage___block_1637_tex;
reg  [5:0] _t___stage___block_1637_vnum0;
reg  [5:0] _t___stage___block_1637_vnum1;
reg  [5:0] _t___stage___block_1637_vnum2;
reg signed [20:0] _t___block_1642_cmp_yx;
reg signed [20:0] _t___block_1642_cmp_zx;
reg signed [20:0] _t___block_1642_cmp_zy;
reg  [0:0] _t___block_1642_x_sel;
reg  [0:0] _t___block_1642_y_sel;
reg  [0:0] _t___block_1642_z_sel;
reg  [5:0] _t___stage___block_1658_tex;
reg  [5:0] _t___stage___block_1658_vnum0;
reg  [5:0] _t___stage___block_1658_vnum1;
reg  [5:0] _t___stage___block_1658_vnum2;
reg signed [20:0] _t___block_1663_cmp_yx;
reg signed [20:0] _t___block_1663_cmp_zx;
reg signed [20:0] _t___block_1663_cmp_zy;
reg  [0:0] _t___block_1663_x_sel;
reg  [0:0] _t___block_1663_y_sel;
reg  [0:0] _t___block_1663_z_sel;
reg  [5:0] _t___stage___block_1679_tex;
reg  [5:0] _t___stage___block_1679_vnum0;
reg  [5:0] _t___stage___block_1679_vnum1;
reg  [5:0] _t___stage___block_1679_vnum2;
reg signed [20:0] _t___block_1684_cmp_yx;
reg signed [20:0] _t___block_1684_cmp_zx;
reg signed [20:0] _t___block_1684_cmp_zy;
reg  [0:0] _t___block_1684_x_sel;
reg  [0:0] _t___block_1684_y_sel;
reg  [0:0] _t___block_1684_z_sel;
reg  [5:0] _t___stage___block_1700_tex;
reg  [5:0] _t___stage___block_1700_vnum0;
reg  [5:0] _t___stage___block_1700_vnum1;
reg  [5:0] _t___stage___block_1700_vnum2;
reg signed [20:0] _t___block_1705_cmp_yx;
reg signed [20:0] _t___block_1705_cmp_zx;
reg signed [20:0] _t___block_1705_cmp_zy;
reg  [0:0] _t___block_1705_x_sel;
reg  [0:0] _t___block_1705_y_sel;
reg  [0:0] _t___block_1705_z_sel;
reg  [5:0] _t___stage___block_1721_tex;
reg  [5:0] _t___stage___block_1721_vnum0;
reg  [5:0] _t___stage___block_1721_vnum1;
reg  [5:0] _t___stage___block_1721_vnum2;
reg signed [20:0] _t___block_1726_cmp_yx;
reg signed [20:0] _t___block_1726_cmp_zx;
reg signed [20:0] _t___block_1726_cmp_zy;
reg  [0:0] _t___block_1726_x_sel;
reg  [0:0] _t___block_1726_y_sel;
reg  [0:0] _t___block_1726_z_sel;
reg  [5:0] _t___stage___block_1742_tex;
reg  [5:0] _t___stage___block_1742_vnum0;
reg  [5:0] _t___stage___block_1742_vnum1;
reg  [5:0] _t___stage___block_1742_vnum2;
reg signed [20:0] _t___block_1747_cmp_yx;
reg signed [20:0] _t___block_1747_cmp_zx;
reg signed [20:0] _t___block_1747_cmp_zy;
reg  [0:0] _t___block_1747_x_sel;
reg  [0:0] _t___block_1747_y_sel;
reg  [0:0] _t___block_1747_z_sel;
reg  [5:0] _t___stage___block_1763_tex;
reg  [5:0] _t___stage___block_1763_vnum0;
reg  [5:0] _t___stage___block_1763_vnum1;
reg  [5:0] _t___stage___block_1763_vnum2;
reg signed [20:0] _t___block_1768_cmp_yx;
reg signed [20:0] _t___block_1768_cmp_zx;
reg signed [20:0] _t___block_1768_cmp_zy;
reg  [0:0] _t___block_1768_x_sel;
reg  [0:0] _t___block_1768_y_sel;
reg  [0:0] _t___block_1768_z_sel;
reg  [5:0] _t___stage___block_1784_tex;
reg  [5:0] _t___stage___block_1784_vnum0;
reg  [5:0] _t___stage___block_1784_vnum1;
reg  [5:0] _t___stage___block_1784_vnum2;
reg signed [20:0] _t___block_1789_cmp_yx;
reg signed [20:0] _t___block_1789_cmp_zx;
reg signed [20:0] _t___block_1789_cmp_zy;
reg  [0:0] _t___block_1789_x_sel;
reg  [0:0] _t___block_1789_y_sel;
reg  [0:0] _t___block_1789_z_sel;
reg  [5:0] _t___stage___block_1805_tex;
reg  [5:0] _t___stage___block_1805_vnum0;
reg  [5:0] _t___stage___block_1805_vnum1;
reg  [5:0] _t___stage___block_1805_vnum2;
reg signed [20:0] _t___block_1810_cmp_yx;
reg signed [20:0] _t___block_1810_cmp_zx;
reg signed [20:0] _t___block_1810_cmp_zy;
reg  [0:0] _t___block_1810_x_sel;
reg  [0:0] _t___block_1810_y_sel;
reg  [0:0] _t___block_1810_z_sel;
reg  [5:0] _t___stage___block_1826_tex;
reg  [5:0] _t___stage___block_1826_vnum0;
reg  [5:0] _t___stage___block_1826_vnum1;
reg  [5:0] _t___stage___block_1826_vnum2;
reg signed [20:0] _t___block_1831_cmp_yx;
reg signed [20:0] _t___block_1831_cmp_zx;
reg signed [20:0] _t___block_1831_cmp_zy;
reg  [0:0] _t___block_1831_x_sel;
reg  [0:0] _t___block_1831_y_sel;
reg  [0:0] _t___block_1831_z_sel;
reg  [5:0] _t___stage___block_1847_tex;
reg  [5:0] _t___stage___block_1847_vnum0;
reg  [5:0] _t___stage___block_1847_vnum1;
reg  [5:0] _t___stage___block_1847_vnum2;
reg signed [20:0] _t___block_1852_cmp_yx;
reg signed [20:0] _t___block_1852_cmp_zx;
reg signed [20:0] _t___block_1852_cmp_zy;
reg  [0:0] _t___block_1852_x_sel;
reg  [0:0] _t___block_1852_y_sel;
reg  [0:0] _t___block_1852_z_sel;
reg  [5:0] _t___stage___block_1868_tex;
reg  [5:0] _t___stage___block_1868_vnum0;
reg  [5:0] _t___stage___block_1868_vnum1;
reg  [5:0] _t___stage___block_1868_vnum2;
reg signed [20:0] _t___block_1873_cmp_yx;
reg signed [20:0] _t___block_1873_cmp_zx;
reg signed [20:0] _t___block_1873_cmp_zy;
reg  [0:0] _t___block_1873_x_sel;
reg  [0:0] _t___block_1873_y_sel;
reg  [0:0] _t___block_1873_z_sel;
reg  [5:0] _t___stage___block_1889_tex;
reg  [5:0] _t___stage___block_1889_vnum0;
reg  [5:0] _t___stage___block_1889_vnum1;
reg  [5:0] _t___stage___block_1889_vnum2;
reg signed [20:0] _t___block_1894_cmp_yx;
reg signed [20:0] _t___block_1894_cmp_zx;
reg signed [20:0] _t___block_1894_cmp_zy;
reg  [0:0] _t___block_1894_x_sel;
reg  [0:0] _t___block_1894_y_sel;
reg  [0:0] _t___block_1894_z_sel;
reg  [5:0] _t___stage___block_1910_tex;
reg  [5:0] _t___stage___block_1910_vnum0;
reg  [5:0] _t___stage___block_1910_vnum1;
reg  [5:0] _t___stage___block_1910_vnum2;
reg signed [20:0] _t___block_1915_cmp_yx;
reg signed [20:0] _t___block_1915_cmp_zx;
reg signed [20:0] _t___block_1915_cmp_zy;
reg  [0:0] _t___block_1915_x_sel;
reg  [0:0] _t___block_1915_y_sel;
reg  [0:0] _t___block_1915_z_sel;
reg  [5:0] _t___stage___block_1931_tex;
reg  [5:0] _t___stage___block_1931_vnum0;
reg  [5:0] _t___stage___block_1931_vnum1;
reg  [5:0] _t___stage___block_1931_vnum2;
reg signed [20:0] _t___block_1936_cmp_yx;
reg signed [20:0] _t___block_1936_cmp_zx;
reg signed [20:0] _t___block_1936_cmp_zy;
reg  [0:0] _t___block_1936_x_sel;
reg  [0:0] _t___block_1936_y_sel;
reg  [0:0] _t___block_1936_z_sel;
reg  [5:0] _t___stage___block_1952_tex;
reg  [5:0] _t___stage___block_1952_vnum0;
reg  [5:0] _t___stage___block_1952_vnum1;
reg  [5:0] _t___stage___block_1952_vnum2;
reg signed [20:0] _t___block_1957_cmp_yx;
reg signed [20:0] _t___block_1957_cmp_zx;
reg signed [20:0] _t___block_1957_cmp_zy;
reg  [0:0] _t___block_1957_x_sel;
reg  [0:0] _t___block_1957_y_sel;
reg  [0:0] _t___block_1957_z_sel;
reg  [5:0] _t___stage___block_1973_tex;
reg  [5:0] _t___stage___block_1973_vnum0;
reg  [5:0] _t___stage___block_1973_vnum1;
reg  [5:0] _t___stage___block_1973_vnum2;
reg signed [20:0] _t___block_1978_cmp_yx;
reg signed [20:0] _t___block_1978_cmp_zx;
reg signed [20:0] _t___block_1978_cmp_zy;
reg  [0:0] _t___block_1978_x_sel;
reg  [0:0] _t___block_1978_y_sel;
reg  [0:0] _t___block_1978_z_sel;
reg  [5:0] _t___stage___block_1994_tex;
reg  [5:0] _t___stage___block_1994_vnum0;
reg  [5:0] _t___stage___block_1994_vnum1;
reg  [5:0] _t___stage___block_1994_vnum2;
reg signed [20:0] _t___block_1999_cmp_yx;
reg signed [20:0] _t___block_1999_cmp_zx;
reg signed [20:0] _t___block_1999_cmp_zy;
reg  [0:0] _t___block_1999_x_sel;
reg  [0:0] _t___block_1999_y_sel;
reg  [0:0] _t___block_1999_z_sel;
reg  [5:0] _t___stage___block_2015_tex;
reg  [5:0] _t___stage___block_2015_vnum0;
reg  [5:0] _t___stage___block_2015_vnum1;
reg  [5:0] _t___stage___block_2015_vnum2;
reg signed [20:0] _t___block_2020_cmp_yx;
reg signed [20:0] _t___block_2020_cmp_zx;
reg signed [20:0] _t___block_2020_cmp_zy;
reg  [0:0] _t___block_2020_x_sel;
reg  [0:0] _t___block_2020_y_sel;
reg  [0:0] _t___block_2020_z_sel;
reg  [5:0] _t___stage___block_2036_tex;
reg  [5:0] _t___stage___block_2036_vnum0;
reg  [5:0] _t___stage___block_2036_vnum1;
reg  [5:0] _t___stage___block_2036_vnum2;
reg signed [20:0] _t___block_2041_cmp_yx;
reg signed [20:0] _t___block_2041_cmp_zx;
reg signed [20:0] _t___block_2041_cmp_zy;
reg  [0:0] _t___block_2041_x_sel;
reg  [0:0] _t___block_2041_y_sel;
reg  [0:0] _t___block_2041_z_sel;
reg  [5:0] _t___stage___block_2057_tex;
reg  [5:0] _t___stage___block_2057_vnum0;
reg  [5:0] _t___stage___block_2057_vnum1;
reg  [5:0] _t___stage___block_2057_vnum2;
reg signed [20:0] _t___block_2062_cmp_yx;
reg signed [20:0] _t___block_2062_cmp_zx;
reg signed [20:0] _t___block_2062_cmp_zy;
reg  [0:0] _t___block_2062_x_sel;
reg  [0:0] _t___block_2062_y_sel;
reg  [0:0] _t___block_2062_z_sel;
reg  [5:0] _t___stage___block_2078_tex;
reg  [5:0] _t___stage___block_2078_vnum0;
reg  [5:0] _t___stage___block_2078_vnum1;
reg  [5:0] _t___stage___block_2078_vnum2;
reg signed [20:0] _t___block_2083_cmp_yx;
reg signed [20:0] _t___block_2083_cmp_zx;
reg signed [20:0] _t___block_2083_cmp_zy;
reg  [0:0] _t___block_2083_x_sel;
reg  [0:0] _t___block_2083_y_sel;
reg  [0:0] _t___block_2083_z_sel;
reg  [5:0] _t___stage___block_2099_tex;
reg  [5:0] _t___stage___block_2099_vnum0;
reg  [5:0] _t___stage___block_2099_vnum1;
reg  [5:0] _t___stage___block_2099_vnum2;
reg signed [20:0] _t___block_2104_cmp_yx;
reg signed [20:0] _t___block_2104_cmp_zx;
reg signed [20:0] _t___block_2104_cmp_zy;
reg  [0:0] _t___block_2104_x_sel;
reg  [0:0] _t___block_2104_y_sel;
reg  [0:0] _t___block_2104_z_sel;
reg  [5:0] _t___stage___block_2120_tex;
reg  [5:0] _t___stage___block_2120_vnum0;
reg  [5:0] _t___stage___block_2120_vnum1;
reg  [5:0] _t___stage___block_2120_vnum2;
reg signed [20:0] _t___block_2125_cmp_yx;
reg signed [20:0] _t___block_2125_cmp_zx;
reg signed [20:0] _t___block_2125_cmp_zy;
reg  [0:0] _t___block_2125_x_sel;
reg  [0:0] _t___block_2125_y_sel;
reg  [0:0] _t___block_2125_z_sel;
reg  [5:0] _t___stage___block_2141_tex;
reg  [5:0] _t___stage___block_2141_vnum0;
reg  [5:0] _t___stage___block_2141_vnum1;
reg  [5:0] _t___stage___block_2141_vnum2;
reg signed [20:0] _t___block_2146_cmp_yx;
reg signed [20:0] _t___block_2146_cmp_zx;
reg signed [20:0] _t___block_2146_cmp_zy;
reg  [0:0] _t___block_2146_x_sel;
reg  [0:0] _t___block_2146_y_sel;
reg  [0:0] _t___block_2146_z_sel;
reg  [5:0] _t___stage___block_2162_tex;
reg  [5:0] _t___stage___block_2162_vnum0;
reg  [5:0] _t___stage___block_2162_vnum1;
reg  [5:0] _t___stage___block_2162_vnum2;
reg signed [20:0] _t___block_2167_cmp_yx;
reg signed [20:0] _t___block_2167_cmp_zx;
reg signed [20:0] _t___block_2167_cmp_zy;
reg  [0:0] _t___block_2167_x_sel;
reg  [0:0] _t___block_2167_y_sel;
reg  [0:0] _t___block_2167_z_sel;
reg  [5:0] _t___stage___block_2183_tex;
reg  [5:0] _t___stage___block_2183_vnum0;
reg  [5:0] _t___stage___block_2183_vnum1;
reg  [5:0] _t___stage___block_2183_vnum2;
reg signed [20:0] _t___block_2188_cmp_yx;
reg signed [20:0] _t___block_2188_cmp_zx;
reg signed [20:0] _t___block_2188_cmp_zy;
reg  [0:0] _t___block_2188_x_sel;
reg  [0:0] _t___block_2188_y_sel;
reg  [0:0] _t___block_2188_z_sel;
reg  [5:0] _t___stage___block_2204_tex;
reg  [5:0] _t___stage___block_2204_vnum0;
reg  [5:0] _t___stage___block_2204_vnum1;
reg  [5:0] _t___stage___block_2204_vnum2;
reg signed [20:0] _t___block_2209_cmp_yx;
reg signed [20:0] _t___block_2209_cmp_zx;
reg signed [20:0] _t___block_2209_cmp_zy;
reg  [0:0] _t___block_2209_x_sel;
reg  [0:0] _t___block_2209_y_sel;
reg  [0:0] _t___block_2209_z_sel;
reg  [5:0] _t___stage___block_2225_tex;
reg  [5:0] _t___stage___block_2225_vnum0;
reg  [5:0] _t___stage___block_2225_vnum1;
reg  [5:0] _t___stage___block_2225_vnum2;
reg signed [20:0] _t___block_2230_cmp_yx;
reg signed [20:0] _t___block_2230_cmp_zx;
reg signed [20:0] _t___block_2230_cmp_zy;
reg  [0:0] _t___block_2230_x_sel;
reg  [0:0] _t___block_2230_y_sel;
reg  [0:0] _t___block_2230_z_sel;
reg  [5:0] _t___stage___block_2246_tex;
reg  [5:0] _t___stage___block_2246_vnum0;
reg  [5:0] _t___stage___block_2246_vnum1;
reg  [5:0] _t___stage___block_2246_vnum2;
reg signed [20:0] _t___block_2251_cmp_yx;
reg signed [20:0] _t___block_2251_cmp_zx;
reg signed [20:0] _t___block_2251_cmp_zy;
reg  [0:0] _t___block_2251_x_sel;
reg  [0:0] _t___block_2251_y_sel;
reg  [0:0] _t___block_2251_z_sel;
reg  [5:0] _t___stage___block_2267_tex;
reg  [5:0] _t___stage___block_2267_vnum0;
reg  [5:0] _t___stage___block_2267_vnum1;
reg  [5:0] _t___stage___block_2267_vnum2;
reg signed [20:0] _t___block_2272_cmp_yx;
reg signed [20:0] _t___block_2272_cmp_zx;
reg signed [20:0] _t___block_2272_cmp_zy;
reg  [0:0] _t___block_2272_x_sel;
reg  [0:0] _t___block_2272_y_sel;
reg  [0:0] _t___block_2272_z_sel;
reg  [5:0] _t___stage___block_2288_tex;
reg  [5:0] _t___stage___block_2288_vnum0;
reg  [5:0] _t___stage___block_2288_vnum1;
reg  [5:0] _t___stage___block_2288_vnum2;
reg signed [20:0] _t___block_2293_cmp_yx;
reg signed [20:0] _t___block_2293_cmp_zx;
reg signed [20:0] _t___block_2293_cmp_zy;
reg  [0:0] _t___block_2293_x_sel;
reg  [0:0] _t___block_2293_y_sel;
reg  [0:0] _t___block_2293_z_sel;
reg  [5:0] _t___stage___block_2309_tex;
reg  [5:0] _t___stage___block_2309_vnum0;
reg  [5:0] _t___stage___block_2309_vnum1;
reg  [5:0] _t___stage___block_2309_vnum2;
reg signed [20:0] _t___block_2314_cmp_yx;
reg signed [20:0] _t___block_2314_cmp_zx;
reg signed [20:0] _t___block_2314_cmp_zy;
reg  [0:0] _t___block_2314_x_sel;
reg  [0:0] _t___block_2314_y_sel;
reg  [0:0] _t___block_2314_z_sel;
reg  [5:0] _t___stage___block_2330_tex;
reg  [5:0] _t___stage___block_2330_vnum0;
reg  [5:0] _t___stage___block_2330_vnum1;
reg  [5:0] _t___stage___block_2330_vnum2;
reg signed [20:0] _t___block_2335_cmp_yx;
reg signed [20:0] _t___block_2335_cmp_zx;
reg signed [20:0] _t___block_2335_cmp_zy;
reg  [0:0] _t___block_2335_x_sel;
reg  [0:0] _t___block_2335_y_sel;
reg  [0:0] _t___block_2335_z_sel;
reg  [5:0] _t___stage___block_2351_tex;
reg  [5:0] _t___stage___block_2351_vnum0;
reg  [5:0] _t___stage___block_2351_vnum1;
reg  [5:0] _t___stage___block_2351_vnum2;
reg signed [20:0] _t___block_2356_cmp_yx;
reg signed [20:0] _t___block_2356_cmp_zx;
reg signed [20:0] _t___block_2356_cmp_zy;
reg  [0:0] _t___block_2356_x_sel;
reg  [0:0] _t___block_2356_y_sel;
reg  [0:0] _t___block_2356_z_sel;
reg  [5:0] _t___stage___block_2372_tex;
reg  [5:0] _t___stage___block_2372_vnum0;
reg  [5:0] _t___stage___block_2372_vnum1;
reg  [5:0] _t___stage___block_2372_vnum2;
reg signed [20:0] _t___block_2377_cmp_yx;
reg signed [20:0] _t___block_2377_cmp_zx;
reg signed [20:0] _t___block_2377_cmp_zy;
reg  [0:0] _t___block_2377_x_sel;
reg  [0:0] _t___block_2377_y_sel;
reg  [0:0] _t___block_2377_z_sel;
reg  [5:0] _t___stage___block_2393_tex;
reg  [5:0] _t___stage___block_2393_vnum0;
reg  [5:0] _t___stage___block_2393_vnum1;
reg  [5:0] _t___stage___block_2393_vnum2;
reg signed [20:0] _t___block_2398_cmp_yx;
reg signed [20:0] _t___block_2398_cmp_zx;
reg signed [20:0] _t___block_2398_cmp_zy;
reg  [0:0] _t___block_2398_x_sel;
reg  [0:0] _t___block_2398_y_sel;
reg  [0:0] _t___block_2398_z_sel;
reg  [5:0] _t___stage___block_2414_tex;
reg  [5:0] _t___stage___block_2414_vnum0;
reg  [5:0] _t___stage___block_2414_vnum1;
reg  [5:0] _t___stage___block_2414_vnum2;
reg signed [20:0] _t___block_2419_cmp_yx;
reg signed [20:0] _t___block_2419_cmp_zx;
reg signed [20:0] _t___block_2419_cmp_zy;
reg  [0:0] _t___block_2419_x_sel;
reg  [0:0] _t___block_2419_y_sel;
reg  [0:0] _t___block_2419_z_sel;
reg  [5:0] _t___stage___block_2435_tex;
reg  [5:0] _t___stage___block_2435_vnum0;
reg  [5:0] _t___stage___block_2435_vnum1;
reg  [5:0] _t___stage___block_2435_vnum2;
reg signed [20:0] _t___block_2440_cmp_yx;
reg signed [20:0] _t___block_2440_cmp_zx;
reg signed [20:0] _t___block_2440_cmp_zy;
reg  [0:0] _t___block_2440_x_sel;
reg  [0:0] _t___block_2440_y_sel;
reg  [0:0] _t___block_2440_z_sel;
reg  [5:0] _t___stage___block_2456_tex;
reg  [5:0] _t___stage___block_2456_vnum0;
reg  [5:0] _t___stage___block_2456_vnum1;
reg  [5:0] _t___stage___block_2456_vnum2;
reg signed [20:0] _t___block_2461_cmp_yx;
reg signed [20:0] _t___block_2461_cmp_zx;
reg signed [20:0] _t___block_2461_cmp_zy;
reg  [0:0] _t___block_2461_x_sel;
reg  [0:0] _t___block_2461_y_sel;
reg  [0:0] _t___block_2461_z_sel;
reg  [5:0] _t___stage___block_2477_tex;
reg  [5:0] _t___stage___block_2477_vnum0;
reg  [5:0] _t___stage___block_2477_vnum1;
reg  [5:0] _t___stage___block_2477_vnum2;
reg signed [20:0] _t___block_2482_cmp_yx;
reg signed [20:0] _t___block_2482_cmp_zx;
reg signed [20:0] _t___block_2482_cmp_zy;
reg  [0:0] _t___block_2482_x_sel;
reg  [0:0] _t___block_2482_y_sel;
reg  [0:0] _t___block_2482_z_sel;
reg  [5:0] _t___stage___block_2498_tex;
reg  [5:0] _t___stage___block_2498_vnum0;
reg  [5:0] _t___stage___block_2498_vnum1;
reg  [5:0] _t___stage___block_2498_vnum2;
reg signed [20:0] _t___block_2503_cmp_yx;
reg signed [20:0] _t___block_2503_cmp_zx;
reg signed [20:0] _t___block_2503_cmp_zy;
reg  [0:0] _t___block_2503_x_sel;
reg  [0:0] _t___block_2503_y_sel;
reg  [0:0] _t___block_2503_z_sel;
reg  [5:0] _t___stage___block_2519_tex;
reg  [5:0] _t___stage___block_2519_vnum0;
reg  [5:0] _t___stage___block_2519_vnum1;
reg  [5:0] _t___stage___block_2519_vnum2;
reg signed [20:0] _t___block_2524_cmp_yx;
reg signed [20:0] _t___block_2524_cmp_zx;
reg signed [20:0] _t___block_2524_cmp_zy;
reg  [0:0] _t___block_2524_x_sel;
reg  [0:0] _t___block_2524_y_sel;
reg  [0:0] _t___block_2524_z_sel;
reg  [5:0] _t___stage___block_2540_tex;
reg  [5:0] _t___stage___block_2540_vnum0;
reg  [5:0] _t___stage___block_2540_vnum1;
reg  [5:0] _t___stage___block_2540_vnum2;
reg signed [20:0] _t___block_2545_cmp_yx;
reg signed [20:0] _t___block_2545_cmp_zx;
reg signed [20:0] _t___block_2545_cmp_zy;
reg  [0:0] _t___block_2545_x_sel;
reg  [0:0] _t___block_2545_y_sel;
reg  [0:0] _t___block_2545_z_sel;
reg  [5:0] _t___stage___block_2561_tex;
reg  [5:0] _t___stage___block_2561_vnum0;
reg  [5:0] _t___stage___block_2561_vnum1;
reg  [5:0] _t___stage___block_2561_vnum2;
reg signed [20:0] _t___block_2566_cmp_yx;
reg signed [20:0] _t___block_2566_cmp_zx;
reg signed [20:0] _t___block_2566_cmp_zy;
reg  [0:0] _t___block_2566_x_sel;
reg  [0:0] _t___block_2566_y_sel;
reg  [0:0] _t___block_2566_z_sel;
reg  [5:0] _t___stage___block_2582_tex;
reg  [5:0] _t___stage___block_2582_vnum0;
reg  [5:0] _t___stage___block_2582_vnum1;
reg  [5:0] _t___stage___block_2582_vnum2;
reg signed [20:0] _t___block_2587_cmp_yx;
reg signed [20:0] _t___block_2587_cmp_zx;
reg signed [20:0] _t___block_2587_cmp_zy;
reg  [0:0] _t___block_2587_x_sel;
reg  [0:0] _t___block_2587_y_sel;
reg  [0:0] _t___block_2587_z_sel;
reg  [5:0] _t___stage___block_2603_tex;
reg  [5:0] _t___stage___block_2603_vnum0;
reg  [5:0] _t___stage___block_2603_vnum1;
reg  [5:0] _t___stage___block_2603_vnum2;
reg signed [20:0] _t___block_2608_cmp_yx;
reg signed [20:0] _t___block_2608_cmp_zx;
reg signed [20:0] _t___block_2608_cmp_zy;
reg  [0:0] _t___block_2608_x_sel;
reg  [0:0] _t___block_2608_y_sel;
reg  [0:0] _t___block_2608_z_sel;
reg  [5:0] _t___stage___block_2624_tex;
reg  [5:0] _t___stage___block_2624_vnum0;
reg  [5:0] _t___stage___block_2624_vnum1;
reg  [5:0] _t___stage___block_2624_vnum2;
reg signed [20:0] _t___block_2629_cmp_yx;
reg signed [20:0] _t___block_2629_cmp_zx;
reg signed [20:0] _t___block_2629_cmp_zy;
reg  [0:0] _t___block_2629_x_sel;
reg  [0:0] _t___block_2629_y_sel;
reg  [0:0] _t___block_2629_z_sel;
reg  [5:0] _t___stage___block_2645_tex;
reg  [5:0] _t___stage___block_2645_vnum0;
reg  [5:0] _t___stage___block_2645_vnum1;
reg  [5:0] _t___stage___block_2645_vnum2;
reg signed [20:0] _t___block_2650_cmp_yx;
reg signed [20:0] _t___block_2650_cmp_zx;
reg signed [20:0] _t___block_2650_cmp_zy;
reg  [0:0] _t___block_2650_x_sel;
reg  [0:0] _t___block_2650_y_sel;
reg  [0:0] _t___block_2650_z_sel;
reg  [5:0] _t___stage___block_2666_tex;
reg  [5:0] _t___stage___block_2666_vnum0;
reg  [5:0] _t___stage___block_2666_vnum1;
reg  [5:0] _t___stage___block_2666_vnum2;
reg signed [20:0] _t___block_2671_cmp_yx;
reg signed [20:0] _t___block_2671_cmp_zx;
reg signed [20:0] _t___block_2671_cmp_zy;
reg  [0:0] _t___block_2671_x_sel;
reg  [0:0] _t___block_2671_y_sel;
reg  [0:0] _t___block_2671_z_sel;
reg  [5:0] _t___stage___block_2687_tex;
reg  [5:0] _t___stage___block_2687_vnum0;
reg  [5:0] _t___stage___block_2687_vnum1;
reg  [5:0] _t___stage___block_2687_vnum2;
reg signed [20:0] _t___block_2692_cmp_yx;
reg signed [20:0] _t___block_2692_cmp_zx;
reg signed [20:0] _t___block_2692_cmp_zy;
reg  [0:0] _t___block_2692_x_sel;
reg  [0:0] _t___block_2692_y_sel;
reg  [0:0] _t___block_2692_z_sel;
reg  [5:0] _t___stage___block_2708_tex;
reg  [5:0] _t___stage___block_2708_vnum0;
reg  [5:0] _t___stage___block_2708_vnum1;
reg  [5:0] _t___stage___block_2708_vnum2;
reg signed [20:0] _t___block_2713_cmp_yx;
reg signed [20:0] _t___block_2713_cmp_zx;
reg signed [20:0] _t___block_2713_cmp_zy;
reg  [0:0] _t___block_2713_x_sel;
reg  [0:0] _t___block_2713_y_sel;
reg  [0:0] _t___block_2713_z_sel;
reg  [7:0] _t___stage___block_2729_fog;
reg  [7:0] _t___stage___block_2729_light;
reg  [15:0] _t___stage___block_2729_shade;
reg  [7:0] _t___block_2731_clr_r;
reg  [7:0] _t___block_2731_clr_g;
reg  [7:0] _t___block_2731_clr_b;
wire  [63:0] _w_tile;

reg signed [23:0] _d_frame = 200;
reg signed [23:0] _q_frame = 200;
reg  [8:0] _d_cos_addr0 = 0;
reg  [8:0] _q_cos_addr0 = 0;
reg  [8:0] _d_cos_addr1 = 0;
reg  [8:0] _q_cos_addr1 = 0;
reg  [8:0] _d_sin_addr0 = 0;
reg  [8:0] _q_sin_addr0 = 0;
reg  [8:0] _d_sin_addr1 = 0;
reg  [8:0] _q_sin_addr1 = 0;
reg  [10:0] _d_invA_addr0 = 0;
reg  [10:0] _q_invA_addr0 = 0;
reg  [10:0] _d_invA_addr1 = 0;
reg  [10:0] _q_invA_addr1 = 0;
reg  [10:0] _d_invB_addr = 0;
reg  [10:0] _q_invB_addr = 0;
reg signed [23:0] _d___pip_5160_1_3___block_25_r_x_delta;
reg signed [23:0] _q___pip_5160_1_3___block_25_r_x_delta;
reg signed [23:0] _d___pip_5160_1_4___block_25_r_x_delta;
reg signed [23:0] _q___pip_5160_1_4___block_25_r_x_delta;
reg signed [23:0] _d___pip_5160_1_3___block_25_r_z_delta;
reg signed [23:0] _q___pip_5160_1_3___block_25_r_z_delta;
reg signed [23:0] _d___pip_5160_1_4___block_25_r_z_delta;
reg signed [23:0] _q___pip_5160_1_4___block_25_r_z_delta;
reg  [7:0] _d___pip_5160_1_135___block_2731_clr_b;
reg  [7:0] _q___pip_5160_1_135___block_2731_clr_b;
reg  [7:0] _d___pip_5160_1_136___block_2731_clr_b;
reg  [7:0] _q___pip_5160_1_136___block_2731_clr_b;
reg  [7:0] _d___pip_5160_1_135___block_2731_clr_g;
reg  [7:0] _q___pip_5160_1_135___block_2731_clr_g;
reg  [7:0] _d___pip_5160_1_136___block_2731_clr_g;
reg  [7:0] _q___pip_5160_1_136___block_2731_clr_g;
reg  [7:0] _d___pip_5160_1_135___block_2731_clr_r;
reg  [7:0] _q___pip_5160_1_135___block_2731_clr_r;
reg  [7:0] _d___pip_5160_1_136___block_2731_clr_r;
reg  [7:0] _q___pip_5160_1_136___block_2731_clr_r;
reg  [19:0] _d___pip_5160_1_6___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_6___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_7___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_7___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_8___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_8___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_9___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_9___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_10___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_10___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_11___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_11___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_12___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_12___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_13___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_13___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_14___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_14___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_15___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_15___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_16___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_16___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_17___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_17___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_18___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_18___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_19___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_19___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_20___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_20___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_21___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_21___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_22___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_22___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_23___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_23___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_24___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_24___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_25___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_25___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_26___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_26___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_27___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_27___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_28___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_28___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_29___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_29___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_30___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_30___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_31___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_31___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_32___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_32___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_33___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_33___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_34___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_34___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_35___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_35___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_36___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_36___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_37___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_37___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_38___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_38___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_39___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_39___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_40___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_40___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_41___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_41___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_42___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_42___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_43___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_43___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_44___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_44___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_45___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_45___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_46___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_46___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_47___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_47___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_48___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_48___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_49___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_49___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_50___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_50___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_51___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_51___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_52___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_52___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_53___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_53___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_54___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_54___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_55___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_55___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_56___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_56___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_57___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_57___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_58___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_58___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_59___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_59___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_60___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_60___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_61___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_61___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_62___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_62___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_63___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_63___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_64___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_64___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_65___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_65___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_66___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_66___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_67___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_67___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_68___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_68___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_69___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_69___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_70___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_70___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_71___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_71___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_72___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_72___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_73___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_73___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_74___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_74___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_75___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_75___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_76___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_76___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_77___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_77___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_78___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_78___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_79___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_79___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_80___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_80___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_81___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_81___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_82___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_82___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_83___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_83___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_84___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_84___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_85___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_85___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_86___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_86___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_87___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_87___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_88___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_88___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_89___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_89___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_90___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_90___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_91___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_91___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_92___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_92___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_93___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_93___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_94___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_94___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_95___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_95___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_96___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_96___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_97___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_97___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_98___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_98___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_99___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_99___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_100___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_100___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_101___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_101___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_102___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_102___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_103___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_103___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_104___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_104___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_105___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_105___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_106___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_106___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_107___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_107___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_108___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_108___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_109___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_109___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_110___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_110___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_111___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_111___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_112___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_112___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_113___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_113___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_114___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_114___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_115___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_115___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_116___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_116___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_117___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_117___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_118___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_118___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_119___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_119___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_120___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_120___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_121___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_121___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_122___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_122___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_123___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_123___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_124___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_124___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_125___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_125___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_126___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_126___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_127___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_127___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_128___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_128___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_129___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_129___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_130___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_130___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_131___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_131___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_132___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_132___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_133___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_133___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_134___block_34_tm_x;
reg  [19:0] _q___pip_5160_1_134___block_34_tm_x;
reg  [19:0] _d___pip_5160_1_6___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_6___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_7___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_7___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_8___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_8___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_9___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_9___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_10___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_10___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_11___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_11___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_12___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_12___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_13___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_13___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_14___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_14___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_15___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_15___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_16___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_16___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_17___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_17___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_18___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_18___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_19___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_19___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_20___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_20___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_21___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_21___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_22___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_22___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_23___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_23___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_24___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_24___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_25___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_25___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_26___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_26___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_27___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_27___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_28___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_28___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_29___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_29___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_30___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_30___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_31___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_31___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_32___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_32___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_33___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_33___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_34___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_34___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_35___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_35___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_36___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_36___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_37___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_37___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_38___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_38___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_39___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_39___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_40___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_40___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_41___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_41___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_42___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_42___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_43___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_43___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_44___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_44___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_45___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_45___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_46___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_46___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_47___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_47___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_48___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_48___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_49___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_49___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_50___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_50___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_51___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_51___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_52___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_52___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_53___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_53___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_54___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_54___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_55___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_55___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_56___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_56___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_57___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_57___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_58___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_58___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_59___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_59___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_60___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_60___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_61___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_61___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_62___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_62___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_63___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_63___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_64___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_64___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_65___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_65___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_66___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_66___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_67___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_67___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_68___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_68___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_69___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_69___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_70___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_70___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_71___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_71___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_72___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_72___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_73___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_73___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_74___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_74___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_75___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_75___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_76___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_76___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_77___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_77___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_78___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_78___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_79___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_79___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_80___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_80___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_81___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_81___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_82___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_82___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_83___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_83___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_84___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_84___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_85___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_85___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_86___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_86___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_87___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_87___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_88___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_88___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_89___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_89___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_90___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_90___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_91___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_91___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_92___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_92___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_93___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_93___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_94___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_94___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_95___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_95___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_96___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_96___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_97___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_97___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_98___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_98___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_99___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_99___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_100___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_100___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_101___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_101___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_102___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_102___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_103___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_103___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_104___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_104___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_105___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_105___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_106___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_106___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_107___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_107___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_108___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_108___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_109___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_109___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_110___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_110___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_111___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_111___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_112___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_112___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_113___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_113___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_114___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_114___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_115___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_115___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_116___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_116___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_117___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_117___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_118___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_118___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_119___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_119___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_120___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_120___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_121___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_121___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_122___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_122___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_123___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_123___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_124___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_124___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_125___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_125___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_126___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_126___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_127___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_127___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_128___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_128___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_129___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_129___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_130___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_130___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_131___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_131___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_132___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_132___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_133___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_133___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_134___block_34_tm_y;
reg  [19:0] _q___pip_5160_1_134___block_34_tm_y;
reg  [19:0] _d___pip_5160_1_6___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_6___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_7___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_7___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_8___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_8___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_9___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_9___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_10___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_10___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_11___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_11___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_12___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_12___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_13___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_13___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_14___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_14___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_15___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_15___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_16___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_16___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_17___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_17___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_18___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_18___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_19___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_19___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_20___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_20___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_21___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_21___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_22___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_22___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_23___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_23___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_24___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_24___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_25___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_25___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_26___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_26___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_27___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_27___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_28___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_28___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_29___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_29___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_30___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_30___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_31___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_31___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_32___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_32___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_33___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_33___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_34___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_34___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_35___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_35___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_36___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_36___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_37___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_37___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_38___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_38___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_39___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_39___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_40___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_40___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_41___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_41___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_42___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_42___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_43___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_43___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_44___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_44___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_45___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_45___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_46___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_46___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_47___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_47___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_48___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_48___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_49___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_49___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_50___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_50___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_51___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_51___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_52___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_52___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_53___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_53___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_54___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_54___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_55___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_55___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_56___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_56___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_57___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_57___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_58___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_58___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_59___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_59___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_60___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_60___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_61___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_61___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_62___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_62___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_63___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_63___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_64___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_64___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_65___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_65___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_66___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_66___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_67___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_67___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_68___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_68___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_69___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_69___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_70___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_70___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_71___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_71___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_72___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_72___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_73___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_73___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_74___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_74___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_75___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_75___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_76___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_76___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_77___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_77___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_78___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_78___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_79___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_79___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_80___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_80___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_81___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_81___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_82___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_82___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_83___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_83___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_84___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_84___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_85___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_85___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_86___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_86___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_87___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_87___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_88___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_88___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_89___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_89___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_90___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_90___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_91___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_91___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_92___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_92___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_93___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_93___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_94___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_94___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_95___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_95___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_96___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_96___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_97___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_97___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_98___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_98___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_99___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_99___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_100___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_100___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_101___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_101___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_102___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_102___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_103___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_103___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_104___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_104___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_105___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_105___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_106___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_106___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_107___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_107___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_108___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_108___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_109___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_109___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_110___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_110___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_111___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_111___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_112___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_112___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_113___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_113___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_114___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_114___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_115___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_115___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_116___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_116___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_117___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_117___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_118___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_118___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_119___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_119___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_120___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_120___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_121___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_121___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_122___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_122___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_123___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_123___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_124___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_124___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_125___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_125___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_126___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_126___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_127___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_127___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_128___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_128___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_129___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_129___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_130___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_130___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_131___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_131___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_132___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_132___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_133___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_133___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_134___block_34_tm_z;
reg  [19:0] _q___pip_5160_1_134___block_34_tm_z;
reg  [19:0] _d___pip_5160_1_6___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_6___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_7___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_7___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_8___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_8___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_9___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_9___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_10___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_10___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_11___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_11___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_12___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_12___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_13___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_13___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_14___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_14___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_15___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_15___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_16___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_16___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_17___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_17___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_18___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_18___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_19___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_19___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_20___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_20___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_21___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_21___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_22___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_22___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_23___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_23___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_24___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_24___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_25___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_25___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_26___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_26___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_27___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_27___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_28___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_28___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_29___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_29___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_30___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_30___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_31___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_31___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_32___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_32___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_33___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_33___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_34___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_34___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_35___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_35___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_36___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_36___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_37___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_37___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_38___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_38___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_39___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_39___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_40___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_40___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_41___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_41___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_42___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_42___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_43___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_43___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_44___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_44___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_45___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_45___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_46___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_46___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_47___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_47___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_48___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_48___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_49___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_49___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_50___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_50___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_51___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_51___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_52___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_52___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_53___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_53___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_54___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_54___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_55___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_55___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_56___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_56___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_57___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_57___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_58___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_58___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_59___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_59___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_60___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_60___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_61___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_61___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_62___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_62___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_63___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_63___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_64___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_64___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_65___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_65___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_66___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_66___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_67___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_67___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_68___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_68___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_69___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_69___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_70___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_70___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_71___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_71___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_72___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_72___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_73___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_73___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_74___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_74___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_75___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_75___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_76___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_76___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_77___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_77___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_78___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_78___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_79___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_79___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_80___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_80___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_81___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_81___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_82___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_82___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_83___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_83___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_84___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_84___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_85___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_85___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_86___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_86___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_87___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_87___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_88___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_88___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_89___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_89___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_90___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_90___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_91___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_91___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_92___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_92___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_93___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_93___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_94___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_94___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_95___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_95___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_96___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_96___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_97___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_97___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_98___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_98___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_99___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_99___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_100___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_100___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_101___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_101___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_102___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_102___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_103___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_103___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_104___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_104___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_105___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_105___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_106___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_106___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_107___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_107___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_108___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_108___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_109___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_109___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_110___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_110___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_111___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_111___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_112___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_112___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_113___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_113___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_114___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_114___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_115___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_115___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_116___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_116___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_117___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_117___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_118___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_118___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_119___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_119___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_120___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_120___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_121___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_121___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_122___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_122___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_123___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_123___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_124___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_124___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_125___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_125___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_126___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_126___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_127___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_127___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_128___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_128___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_129___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_129___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_130___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_130___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_131___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_131___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_132___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_132___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_133___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_133___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_134___block_40_dt_x;
reg  [19:0] _q___pip_5160_1_134___block_40_dt_x;
reg  [19:0] _d___pip_5160_1_6___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_6___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_7___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_7___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_8___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_8___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_9___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_9___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_10___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_10___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_11___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_11___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_12___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_12___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_13___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_13___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_14___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_14___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_15___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_15___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_16___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_16___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_17___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_17___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_18___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_18___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_19___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_19___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_20___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_20___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_21___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_21___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_22___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_22___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_23___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_23___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_24___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_24___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_25___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_25___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_26___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_26___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_27___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_27___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_28___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_28___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_29___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_29___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_30___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_30___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_31___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_31___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_32___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_32___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_33___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_33___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_34___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_34___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_35___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_35___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_36___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_36___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_37___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_37___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_38___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_38___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_39___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_39___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_40___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_40___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_41___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_41___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_42___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_42___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_43___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_43___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_44___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_44___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_45___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_45___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_46___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_46___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_47___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_47___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_48___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_48___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_49___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_49___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_50___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_50___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_51___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_51___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_52___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_52___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_53___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_53___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_54___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_54___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_55___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_55___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_56___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_56___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_57___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_57___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_58___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_58___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_59___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_59___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_60___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_60___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_61___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_61___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_62___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_62___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_63___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_63___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_64___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_64___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_65___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_65___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_66___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_66___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_67___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_67___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_68___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_68___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_69___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_69___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_70___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_70___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_71___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_71___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_72___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_72___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_73___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_73___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_74___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_74___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_75___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_75___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_76___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_76___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_77___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_77___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_78___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_78___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_79___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_79___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_80___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_80___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_81___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_81___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_82___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_82___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_83___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_83___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_84___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_84___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_85___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_85___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_86___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_86___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_87___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_87___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_88___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_88___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_89___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_89___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_90___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_90___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_91___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_91___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_92___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_92___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_93___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_93___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_94___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_94___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_95___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_95___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_96___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_96___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_97___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_97___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_98___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_98___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_99___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_99___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_100___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_100___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_101___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_101___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_102___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_102___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_103___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_103___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_104___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_104___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_105___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_105___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_106___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_106___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_107___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_107___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_108___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_108___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_109___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_109___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_110___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_110___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_111___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_111___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_112___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_112___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_113___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_113___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_114___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_114___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_115___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_115___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_116___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_116___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_117___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_117___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_118___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_118___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_119___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_119___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_120___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_120___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_121___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_121___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_122___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_122___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_123___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_123___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_124___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_124___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_125___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_125___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_126___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_126___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_127___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_127___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_128___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_128___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_129___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_129___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_130___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_130___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_131___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_131___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_132___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_132___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_133___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_133___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_134___block_40_dt_y;
reg  [19:0] _q___pip_5160_1_134___block_40_dt_y;
reg  [19:0] _d___pip_5160_1_6___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_6___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_7___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_7___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_8___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_8___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_9___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_9___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_10___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_10___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_11___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_11___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_12___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_12___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_13___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_13___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_14___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_14___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_15___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_15___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_16___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_16___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_17___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_17___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_18___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_18___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_19___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_19___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_20___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_20___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_21___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_21___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_22___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_22___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_23___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_23___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_24___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_24___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_25___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_25___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_26___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_26___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_27___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_27___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_28___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_28___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_29___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_29___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_30___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_30___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_31___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_31___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_32___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_32___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_33___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_33___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_34___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_34___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_35___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_35___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_36___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_36___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_37___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_37___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_38___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_38___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_39___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_39___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_40___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_40___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_41___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_41___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_42___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_42___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_43___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_43___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_44___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_44___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_45___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_45___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_46___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_46___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_47___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_47___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_48___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_48___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_49___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_49___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_50___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_50___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_51___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_51___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_52___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_52___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_53___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_53___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_54___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_54___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_55___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_55___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_56___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_56___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_57___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_57___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_58___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_58___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_59___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_59___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_60___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_60___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_61___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_61___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_62___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_62___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_63___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_63___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_64___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_64___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_65___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_65___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_66___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_66___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_67___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_67___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_68___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_68___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_69___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_69___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_70___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_70___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_71___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_71___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_72___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_72___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_73___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_73___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_74___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_74___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_75___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_75___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_76___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_76___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_77___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_77___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_78___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_78___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_79___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_79___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_80___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_80___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_81___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_81___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_82___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_82___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_83___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_83___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_84___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_84___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_85___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_85___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_86___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_86___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_87___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_87___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_88___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_88___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_89___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_89___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_90___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_90___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_91___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_91___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_92___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_92___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_93___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_93___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_94___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_94___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_95___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_95___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_96___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_96___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_97___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_97___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_98___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_98___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_99___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_99___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_100___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_100___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_101___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_101___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_102___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_102___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_103___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_103___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_104___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_104___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_105___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_105___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_106___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_106___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_107___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_107___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_108___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_108___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_109___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_109___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_110___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_110___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_111___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_111___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_112___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_112___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_113___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_113___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_114___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_114___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_115___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_115___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_116___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_116___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_117___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_117___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_118___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_118___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_119___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_119___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_120___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_120___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_121___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_121___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_122___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_122___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_123___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_123___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_124___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_124___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_125___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_125___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_126___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_126___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_127___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_127___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_128___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_128___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_129___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_129___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_130___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_130___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_131___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_131___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_132___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_132___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_133___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_133___block_40_dt_z;
reg  [19:0] _d___pip_5160_1_134___block_40_dt_z;
reg  [19:0] _q___pip_5160_1_134___block_40_dt_z;
reg  [13:0] _d___pip_5160_1_4___stage___block_26_brd_x;
reg  [13:0] _q___pip_5160_1_4___stage___block_26_brd_x;
reg  [13:0] _d___pip_5160_1_5___stage___block_26_brd_x;
reg  [13:0] _q___pip_5160_1_5___stage___block_26_brd_x;
reg  [13:0] _d___pip_5160_1_6___stage___block_26_brd_x;
reg  [13:0] _q___pip_5160_1_6___stage___block_26_brd_x;
reg  [13:0] _d___pip_5160_1_4___stage___block_26_brd_y;
reg  [13:0] _q___pip_5160_1_4___stage___block_26_brd_y;
reg  [13:0] _d___pip_5160_1_5___stage___block_26_brd_y;
reg  [13:0] _q___pip_5160_1_5___stage___block_26_brd_y;
reg  [13:0] _d___pip_5160_1_6___stage___block_26_brd_y;
reg  [13:0] _q___pip_5160_1_6___stage___block_26_brd_y;
reg  [13:0] _d___pip_5160_1_4___stage___block_26_brd_z;
reg  [13:0] _q___pip_5160_1_4___stage___block_26_brd_z;
reg  [13:0] _d___pip_5160_1_5___stage___block_26_brd_z;
reg  [13:0] _q___pip_5160_1_5___stage___block_26_brd_z;
reg  [13:0] _d___pip_5160_1_6___stage___block_26_brd_z;
reg  [13:0] _q___pip_5160_1_6___stage___block_26_brd_z;
reg signed [15:0] _d___pip_5160_1_4___stage___block_26_rd_x;
reg signed [15:0] _q___pip_5160_1_4___stage___block_26_rd_x;
reg signed [15:0] _d___pip_5160_1_5___stage___block_26_rd_x;
reg signed [15:0] _q___pip_5160_1_5___stage___block_26_rd_x;
reg signed [15:0] _d___pip_5160_1_4___stage___block_26_rd_y;
reg signed [15:0] _q___pip_5160_1_4___stage___block_26_rd_y;
reg signed [15:0] _d___pip_5160_1_5___stage___block_26_rd_y;
reg signed [15:0] _q___pip_5160_1_5___stage___block_26_rd_y;
reg signed [15:0] _d___pip_5160_1_4___stage___block_26_rd_z;
reg signed [15:0] _q___pip_5160_1_4___stage___block_26_rd_z;
reg signed [15:0] _d___pip_5160_1_5___stage___block_26_rd_z;
reg signed [15:0] _q___pip_5160_1_5___stage___block_26_rd_z;
reg signed [1:0] _d___pip_5160_1_4___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_4___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_5___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_5___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_6___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_6___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_7___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_7___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_8___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_8___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_9___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_9___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_10___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_10___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_11___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_11___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_12___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_12___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_13___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_13___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_14___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_14___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_15___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_15___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_16___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_16___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_17___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_17___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_18___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_18___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_19___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_19___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_20___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_20___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_21___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_21___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_22___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_22___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_23___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_23___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_24___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_24___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_25___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_25___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_26___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_26___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_27___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_27___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_28___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_28___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_29___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_29___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_30___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_30___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_31___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_31___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_32___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_32___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_33___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_33___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_34___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_34___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_35___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_35___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_36___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_36___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_37___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_37___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_38___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_38___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_39___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_39___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_40___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_40___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_41___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_41___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_42___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_42___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_43___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_43___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_44___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_44___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_45___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_45___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_46___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_46___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_47___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_47___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_48___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_48___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_49___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_49___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_50___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_50___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_51___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_51___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_52___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_52___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_53___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_53___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_54___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_54___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_55___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_55___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_56___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_56___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_57___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_57___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_58___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_58___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_59___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_59___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_60___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_60___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_61___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_61___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_62___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_62___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_63___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_63___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_64___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_64___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_65___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_65___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_66___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_66___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_67___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_67___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_68___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_68___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_69___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_69___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_70___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_70___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_71___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_71___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_72___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_72___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_73___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_73___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_74___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_74___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_75___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_75___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_76___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_76___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_77___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_77___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_78___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_78___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_79___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_79___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_80___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_80___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_81___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_81___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_82___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_82___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_83___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_83___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_84___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_84___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_85___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_85___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_86___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_86___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_87___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_87___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_88___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_88___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_89___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_89___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_90___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_90___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_91___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_91___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_92___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_92___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_93___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_93___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_94___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_94___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_95___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_95___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_96___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_96___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_97___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_97___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_98___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_98___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_99___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_99___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_100___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_100___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_101___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_101___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_102___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_102___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_103___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_103___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_104___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_104___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_105___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_105___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_106___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_106___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_107___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_107___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_108___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_108___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_109___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_109___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_110___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_110___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_111___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_111___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_112___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_112___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_113___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_113___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_114___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_114___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_115___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_115___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_116___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_116___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_117___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_117___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_118___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_118___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_119___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_119___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_120___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_120___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_121___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_121___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_122___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_122___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_123___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_123___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_124___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_124___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_125___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_125___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_126___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_126___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_127___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_127___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_128___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_128___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_129___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_129___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_130___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_130___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_131___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_131___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_132___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_132___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_133___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_133___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_134___stage___block_26_s_x;
reg signed [1:0] _q___pip_5160_1_134___stage___block_26_s_x;
reg signed [1:0] _d___pip_5160_1_4___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_4___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_5___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_5___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_6___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_6___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_7___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_7___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_8___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_8___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_9___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_9___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_10___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_10___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_11___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_11___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_12___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_12___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_13___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_13___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_14___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_14___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_15___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_15___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_16___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_16___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_17___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_17___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_18___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_18___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_19___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_19___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_20___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_20___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_21___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_21___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_22___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_22___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_23___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_23___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_24___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_24___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_25___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_25___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_26___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_26___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_27___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_27___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_28___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_28___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_29___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_29___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_30___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_30___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_31___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_31___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_32___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_32___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_33___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_33___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_34___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_34___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_35___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_35___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_36___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_36___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_37___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_37___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_38___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_38___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_39___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_39___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_40___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_40___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_41___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_41___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_42___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_42___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_43___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_43___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_44___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_44___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_45___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_45___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_46___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_46___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_47___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_47___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_48___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_48___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_49___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_49___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_50___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_50___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_51___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_51___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_52___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_52___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_53___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_53___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_54___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_54___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_55___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_55___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_56___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_56___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_57___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_57___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_58___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_58___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_59___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_59___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_60___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_60___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_61___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_61___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_62___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_62___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_63___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_63___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_64___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_64___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_65___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_65___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_66___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_66___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_67___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_67___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_68___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_68___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_69___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_69___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_70___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_70___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_71___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_71___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_72___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_72___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_73___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_73___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_74___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_74___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_75___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_75___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_76___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_76___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_77___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_77___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_78___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_78___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_79___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_79___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_80___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_80___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_81___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_81___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_82___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_82___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_83___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_83___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_84___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_84___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_85___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_85___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_86___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_86___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_87___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_87___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_88___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_88___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_89___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_89___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_90___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_90___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_91___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_91___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_92___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_92___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_93___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_93___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_94___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_94___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_95___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_95___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_96___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_96___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_97___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_97___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_98___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_98___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_99___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_99___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_100___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_100___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_101___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_101___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_102___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_102___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_103___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_103___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_104___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_104___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_105___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_105___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_106___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_106___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_107___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_107___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_108___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_108___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_109___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_109___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_110___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_110___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_111___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_111___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_112___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_112___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_113___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_113___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_114___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_114___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_115___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_115___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_116___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_116___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_117___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_117___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_118___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_118___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_119___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_119___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_120___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_120___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_121___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_121___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_122___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_122___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_123___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_123___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_124___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_124___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_125___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_125___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_126___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_126___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_127___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_127___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_128___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_128___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_129___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_129___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_130___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_130___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_131___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_131___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_132___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_132___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_133___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_133___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_134___stage___block_26_s_y;
reg signed [1:0] _q___pip_5160_1_134___stage___block_26_s_y;
reg signed [1:0] _d___pip_5160_1_4___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_4___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_5___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_5___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_6___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_6___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_7___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_7___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_8___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_8___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_9___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_9___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_10___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_10___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_11___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_11___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_12___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_12___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_13___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_13___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_14___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_14___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_15___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_15___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_16___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_16___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_17___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_17___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_18___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_18___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_19___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_19___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_20___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_20___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_21___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_21___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_22___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_22___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_23___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_23___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_24___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_24___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_25___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_25___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_26___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_26___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_27___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_27___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_28___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_28___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_29___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_29___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_30___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_30___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_31___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_31___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_32___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_32___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_33___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_33___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_34___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_34___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_35___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_35___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_36___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_36___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_37___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_37___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_38___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_38___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_39___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_39___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_40___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_40___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_41___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_41___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_42___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_42___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_43___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_43___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_44___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_44___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_45___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_45___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_46___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_46___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_47___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_47___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_48___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_48___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_49___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_49___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_50___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_50___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_51___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_51___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_52___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_52___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_53___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_53___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_54___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_54___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_55___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_55___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_56___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_56___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_57___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_57___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_58___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_58___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_59___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_59___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_60___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_60___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_61___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_61___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_62___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_62___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_63___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_63___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_64___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_64___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_65___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_65___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_66___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_66___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_67___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_67___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_68___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_68___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_69___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_69___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_70___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_70___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_71___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_71___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_72___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_72___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_73___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_73___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_74___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_74___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_75___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_75___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_76___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_76___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_77___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_77___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_78___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_78___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_79___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_79___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_80___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_80___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_81___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_81___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_82___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_82___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_83___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_83___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_84___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_84___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_85___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_85___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_86___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_86___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_87___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_87___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_88___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_88___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_89___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_89___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_90___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_90___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_91___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_91___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_92___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_92___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_93___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_93___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_94___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_94___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_95___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_95___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_96___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_96___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_97___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_97___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_98___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_98___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_99___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_99___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_100___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_100___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_101___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_101___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_102___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_102___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_103___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_103___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_104___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_104___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_105___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_105___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_106___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_106___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_107___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_107___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_108___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_108___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_109___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_109___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_110___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_110___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_111___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_111___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_112___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_112___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_113___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_113___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_114___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_114___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_115___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_115___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_116___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_116___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_117___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_117___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_118___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_118___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_119___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_119___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_120___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_120___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_121___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_121___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_122___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_122___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_123___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_123___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_124___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_124___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_125___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_125___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_126___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_126___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_127___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_127___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_128___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_128___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_129___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_129___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_130___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_130___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_131___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_131___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_132___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_132___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_133___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_133___stage___block_26_s_z;
reg signed [1:0] _d___pip_5160_1_134___stage___block_26_s_z;
reg signed [1:0] _q___pip_5160_1_134___stage___block_26_s_z;
reg signed [11:0] _d___pip_5160_1_4___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_4___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_5___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_5___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_6___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_6___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_7___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_7___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_8___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_8___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_9___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_9___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_10___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_10___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_11___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_11___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_12___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_12___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_13___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_13___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_14___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_14___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_15___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_15___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_16___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_16___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_17___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_17___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_18___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_18___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_19___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_19___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_20___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_20___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_21___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_21___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_22___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_22___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_23___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_23___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_24___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_24___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_25___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_25___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_26___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_26___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_27___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_27___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_28___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_28___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_29___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_29___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_30___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_30___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_31___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_31___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_32___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_32___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_33___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_33___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_34___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_34___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_35___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_35___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_36___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_36___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_37___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_37___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_38___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_38___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_39___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_39___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_40___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_40___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_41___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_41___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_42___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_42___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_43___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_43___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_44___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_44___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_45___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_45___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_46___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_46___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_47___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_47___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_48___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_48___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_49___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_49___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_50___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_50___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_51___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_51___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_52___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_52___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_53___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_53___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_54___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_54___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_55___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_55___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_56___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_56___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_57___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_57___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_58___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_58___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_59___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_59___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_60___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_60___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_61___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_61___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_62___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_62___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_63___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_63___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_64___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_64___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_65___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_65___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_66___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_66___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_67___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_67___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_68___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_68___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_69___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_69___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_70___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_70___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_71___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_71___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_72___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_72___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_73___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_73___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_74___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_74___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_75___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_75___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_76___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_76___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_77___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_77___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_78___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_78___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_79___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_79___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_80___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_80___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_81___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_81___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_82___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_82___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_83___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_83___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_84___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_84___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_85___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_85___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_86___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_86___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_87___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_87___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_88___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_88___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_89___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_89___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_90___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_90___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_91___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_91___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_92___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_92___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_93___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_93___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_94___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_94___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_95___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_95___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_96___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_96___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_97___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_97___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_98___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_98___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_99___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_99___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_100___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_100___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_101___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_101___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_102___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_102___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_103___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_103___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_104___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_104___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_105___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_105___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_106___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_106___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_107___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_107___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_108___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_108___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_109___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_109___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_110___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_110___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_111___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_111___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_112___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_112___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_113___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_113___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_114___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_114___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_115___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_115___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_116___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_116___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_117___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_117___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_118___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_118___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_119___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_119___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_120___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_120___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_121___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_121___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_122___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_122___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_123___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_123___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_124___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_124___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_125___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_125___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_126___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_126___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_127___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_127___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_128___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_128___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_129___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_129___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_130___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_130___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_131___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_131___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_132___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_132___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_133___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_133___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_134___stage___block_26_v_x;
reg signed [11:0] _q___pip_5160_1_134___stage___block_26_v_x;
reg signed [11:0] _d___pip_5160_1_4___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_4___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_5___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_5___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_6___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_6___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_7___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_7___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_8___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_8___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_9___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_9___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_10___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_10___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_11___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_11___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_12___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_12___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_13___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_13___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_14___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_14___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_15___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_15___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_16___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_16___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_17___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_17___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_18___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_18___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_19___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_19___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_20___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_20___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_21___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_21___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_22___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_22___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_23___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_23___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_24___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_24___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_25___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_25___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_26___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_26___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_27___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_27___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_28___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_28___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_29___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_29___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_30___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_30___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_31___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_31___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_32___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_32___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_33___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_33___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_34___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_34___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_35___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_35___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_36___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_36___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_37___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_37___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_38___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_38___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_39___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_39___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_40___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_40___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_41___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_41___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_42___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_42___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_43___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_43___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_44___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_44___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_45___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_45___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_46___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_46___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_47___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_47___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_48___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_48___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_49___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_49___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_50___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_50___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_51___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_51___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_52___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_52___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_53___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_53___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_54___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_54___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_55___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_55___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_56___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_56___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_57___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_57___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_58___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_58___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_59___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_59___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_60___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_60___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_61___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_61___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_62___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_62___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_63___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_63___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_64___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_64___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_65___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_65___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_66___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_66___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_67___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_67___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_68___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_68___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_69___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_69___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_70___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_70___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_71___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_71___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_72___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_72___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_73___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_73___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_74___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_74___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_75___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_75___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_76___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_76___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_77___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_77___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_78___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_78___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_79___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_79___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_80___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_80___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_81___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_81___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_82___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_82___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_83___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_83___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_84___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_84___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_85___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_85___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_86___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_86___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_87___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_87___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_88___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_88___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_89___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_89___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_90___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_90___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_91___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_91___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_92___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_92___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_93___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_93___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_94___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_94___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_95___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_95___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_96___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_96___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_97___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_97___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_98___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_98___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_99___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_99___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_100___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_100___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_101___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_101___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_102___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_102___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_103___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_103___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_104___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_104___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_105___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_105___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_106___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_106___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_107___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_107___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_108___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_108___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_109___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_109___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_110___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_110___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_111___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_111___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_112___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_112___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_113___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_113___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_114___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_114___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_115___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_115___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_116___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_116___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_117___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_117___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_118___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_118___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_119___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_119___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_120___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_120___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_121___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_121___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_122___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_122___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_123___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_123___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_124___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_124___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_125___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_125___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_126___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_126___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_127___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_127___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_128___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_128___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_129___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_129___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_130___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_130___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_131___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_131___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_132___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_132___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_133___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_133___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_134___stage___block_26_v_y;
reg signed [11:0] _q___pip_5160_1_134___stage___block_26_v_y;
reg signed [11:0] _d___pip_5160_1_4___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_4___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_5___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_5___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_6___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_6___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_7___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_7___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_8___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_8___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_9___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_9___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_10___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_10___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_11___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_11___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_12___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_12___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_13___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_13___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_14___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_14___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_15___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_15___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_16___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_16___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_17___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_17___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_18___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_18___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_19___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_19___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_20___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_20___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_21___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_21___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_22___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_22___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_23___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_23___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_24___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_24___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_25___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_25___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_26___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_26___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_27___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_27___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_28___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_28___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_29___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_29___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_30___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_30___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_31___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_31___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_32___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_32___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_33___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_33___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_34___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_34___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_35___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_35___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_36___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_36___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_37___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_37___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_38___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_38___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_39___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_39___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_40___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_40___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_41___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_41___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_42___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_42___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_43___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_43___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_44___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_44___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_45___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_45___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_46___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_46___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_47___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_47___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_48___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_48___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_49___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_49___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_50___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_50___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_51___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_51___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_52___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_52___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_53___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_53___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_54___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_54___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_55___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_55___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_56___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_56___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_57___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_57___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_58___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_58___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_59___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_59___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_60___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_60___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_61___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_61___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_62___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_62___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_63___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_63___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_64___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_64___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_65___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_65___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_66___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_66___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_67___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_67___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_68___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_68___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_69___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_69___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_70___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_70___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_71___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_71___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_72___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_72___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_73___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_73___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_74___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_74___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_75___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_75___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_76___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_76___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_77___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_77___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_78___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_78___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_79___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_79___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_80___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_80___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_81___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_81___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_82___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_82___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_83___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_83___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_84___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_84___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_85___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_85___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_86___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_86___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_87___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_87___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_88___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_88___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_89___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_89___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_90___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_90___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_91___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_91___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_92___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_92___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_93___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_93___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_94___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_94___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_95___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_95___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_96___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_96___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_97___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_97___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_98___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_98___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_99___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_99___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_100___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_100___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_101___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_101___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_102___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_102___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_103___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_103___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_104___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_104___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_105___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_105___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_106___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_106___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_107___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_107___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_108___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_108___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_109___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_109___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_110___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_110___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_111___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_111___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_112___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_112___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_113___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_113___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_114___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_114___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_115___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_115___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_116___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_116___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_117___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_117___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_118___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_118___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_119___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_119___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_120___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_120___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_121___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_121___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_122___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_122___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_123___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_123___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_124___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_124___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_125___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_125___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_126___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_126___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_127___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_127___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_128___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_128___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_129___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_129___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_130___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_130___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_131___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_131___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_132___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_132___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_133___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_133___stage___block_26_v_z;
reg signed [11:0] _d___pip_5160_1_134___stage___block_26_v_z;
reg signed [11:0] _q___pip_5160_1_134___stage___block_26_v_z;
reg  [7:0] _d___pip_5160_1_0___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_0___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_1___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_1___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_2___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_2___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_3___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_3___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_4___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_4___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_5___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_5___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_6___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_6___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_7___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_7___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_8___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_8___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_9___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_9___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_10___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_10___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_11___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_11___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_12___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_12___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_13___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_13___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_14___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_14___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_15___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_15___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_16___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_16___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_17___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_17___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_18___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_18___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_19___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_19___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_20___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_20___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_21___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_21___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_22___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_22___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_23___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_23___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_24___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_24___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_25___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_25___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_26___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_26___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_27___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_27___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_28___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_28___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_29___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_29___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_30___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_30___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_31___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_31___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_32___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_32___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_33___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_33___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_34___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_34___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_35___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_35___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_36___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_36___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_37___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_37___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_38___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_38___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_39___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_39___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_40___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_40___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_41___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_41___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_42___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_42___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_43___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_43___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_44___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_44___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_45___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_45___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_46___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_46___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_47___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_47___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_48___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_48___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_49___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_49___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_50___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_50___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_51___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_51___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_52___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_52___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_53___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_53___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_54___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_54___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_55___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_55___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_56___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_56___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_57___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_57___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_58___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_58___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_59___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_59___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_60___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_60___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_61___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_61___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_62___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_62___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_63___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_63___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_64___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_64___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_65___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_65___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_66___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_66___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_67___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_67___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_68___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_68___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_69___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_69___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_70___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_70___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_71___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_71___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_72___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_72___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_73___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_73___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_74___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_74___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_75___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_75___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_76___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_76___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_77___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_77___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_78___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_78___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_79___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_79___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_80___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_80___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_81___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_81___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_82___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_82___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_83___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_83___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_84___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_84___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_85___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_85___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_86___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_86___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_87___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_87___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_88___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_88___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_89___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_89___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_90___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_90___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_91___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_91___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_92___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_92___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_93___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_93___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_94___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_94___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_95___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_95___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_96___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_96___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_97___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_97___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_98___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_98___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_99___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_99___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_100___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_100___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_101___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_101___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_102___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_102___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_103___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_103___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_104___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_104___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_105___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_105___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_106___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_106___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_107___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_107___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_108___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_108___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_109___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_109___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_110___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_110___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_111___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_111___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_112___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_112___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_113___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_113___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_114___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_114___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_115___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_115___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_116___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_116___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_117___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_117___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_118___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_118___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_119___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_119___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_120___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_120___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_121___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_121___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_122___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_122___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_123___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_123___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_124___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_124___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_125___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_125___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_126___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_126___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_127___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_127___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_128___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_128___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_129___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_129___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_130___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_130___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_131___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_131___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_132___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_132___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_133___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_133___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_134___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_134___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_135___stage___block_6_clr;
reg  [7:0] _q___pip_5160_1_135___stage___block_6_clr;
reg  [7:0] _d___pip_5160_1_0___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_0___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_1___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_1___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_2___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_2___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_3___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_3___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_4___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_4___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_5___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_5___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_6___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_6___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_7___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_7___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_8___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_8___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_9___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_9___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_10___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_10___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_11___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_11___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_12___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_12___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_13___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_13___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_14___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_14___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_15___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_15___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_16___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_16___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_17___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_17___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_18___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_18___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_19___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_19___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_20___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_20___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_21___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_21___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_22___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_22___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_23___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_23___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_24___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_24___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_25___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_25___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_26___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_26___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_27___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_27___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_28___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_28___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_29___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_29___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_30___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_30___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_31___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_31___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_32___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_32___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_33___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_33___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_34___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_34___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_35___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_35___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_36___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_36___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_37___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_37___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_38___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_38___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_39___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_39___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_40___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_40___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_41___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_41___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_42___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_42___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_43___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_43___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_44___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_44___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_45___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_45___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_46___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_46___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_47___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_47___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_48___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_48___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_49___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_49___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_50___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_50___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_51___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_51___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_52___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_52___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_53___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_53___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_54___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_54___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_55___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_55___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_56___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_56___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_57___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_57___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_58___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_58___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_59___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_59___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_60___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_60___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_61___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_61___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_62___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_62___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_63___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_63___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_64___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_64___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_65___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_65___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_66___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_66___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_67___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_67___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_68___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_68___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_69___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_69___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_70___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_70___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_71___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_71___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_72___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_72___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_73___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_73___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_74___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_74___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_75___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_75___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_76___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_76___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_77___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_77___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_78___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_78___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_79___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_79___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_80___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_80___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_81___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_81___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_82___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_82___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_83___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_83___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_84___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_84___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_85___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_85___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_86___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_86___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_87___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_87___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_88___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_88___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_89___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_89___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_90___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_90___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_91___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_91___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_92___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_92___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_93___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_93___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_94___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_94___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_95___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_95___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_96___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_96___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_97___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_97___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_98___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_98___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_99___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_99___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_100___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_100___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_101___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_101___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_102___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_102___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_103___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_103___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_104___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_104___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_105___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_105___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_106___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_106___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_107___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_107___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_108___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_108___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_109___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_109___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_110___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_110___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_111___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_111___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_112___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_112___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_113___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_113___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_114___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_114___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_115___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_115___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_116___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_116___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_117___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_117___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_118___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_118___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_119___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_119___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_120___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_120___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_121___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_121___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_122___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_122___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_123___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_123___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_124___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_124___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_125___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_125___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_126___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_126___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_127___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_127___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_128___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_128___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_129___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_129___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_130___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_130___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_131___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_131___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_132___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_132___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_133___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_133___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_134___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_134___stage___block_6_dist;
reg  [7:0] _d___pip_5160_1_135___stage___block_6_dist;
reg  [7:0] _q___pip_5160_1_135___stage___block_6_dist;
reg  [0:0] _d___pip_5160_1_0___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_0___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_1___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_1___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_2___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_2___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_3___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_3___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_4___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_4___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_5___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_5___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_6___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_6___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_7___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_7___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_8___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_8___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_9___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_9___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_10___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_10___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_11___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_11___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_12___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_12___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_13___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_13___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_14___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_14___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_15___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_15___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_16___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_16___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_17___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_17___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_18___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_18___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_19___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_19___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_20___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_20___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_21___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_21___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_22___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_22___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_23___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_23___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_24___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_24___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_25___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_25___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_26___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_26___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_27___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_27___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_28___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_28___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_29___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_29___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_30___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_30___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_31___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_31___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_32___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_32___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_33___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_33___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_34___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_34___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_35___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_35___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_36___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_36___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_37___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_37___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_38___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_38___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_39___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_39___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_40___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_40___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_41___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_41___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_42___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_42___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_43___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_43___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_44___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_44___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_45___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_45___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_46___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_46___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_47___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_47___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_48___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_48___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_49___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_49___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_50___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_50___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_51___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_51___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_52___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_52___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_53___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_53___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_54___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_54___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_55___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_55___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_56___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_56___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_57___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_57___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_58___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_58___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_59___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_59___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_60___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_60___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_61___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_61___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_62___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_62___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_63___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_63___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_64___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_64___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_65___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_65___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_66___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_66___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_67___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_67___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_68___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_68___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_69___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_69___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_70___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_70___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_71___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_71___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_72___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_72___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_73___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_73___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_74___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_74___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_75___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_75___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_76___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_76___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_77___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_77___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_78___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_78___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_79___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_79___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_80___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_80___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_81___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_81___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_82___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_82___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_83___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_83___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_84___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_84___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_85___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_85___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_86___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_86___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_87___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_87___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_88___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_88___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_89___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_89___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_90___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_90___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_91___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_91___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_92___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_92___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_93___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_93___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_94___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_94___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_95___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_95___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_96___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_96___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_97___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_97___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_98___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_98___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_99___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_99___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_100___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_100___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_101___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_101___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_102___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_102___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_103___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_103___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_104___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_104___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_105___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_105___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_106___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_106___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_107___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_107___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_108___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_108___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_109___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_109___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_110___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_110___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_111___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_111___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_112___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_112___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_113___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_113___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_114___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_114___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_115___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_115___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_116___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_116___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_117___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_117___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_118___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_118___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_119___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_119___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_120___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_120___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_121___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_121___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_122___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_122___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_123___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_123___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_124___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_124___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_125___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_125___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_126___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_126___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_127___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_127___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_128___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_128___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_129___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_129___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_130___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_130___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_131___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_131___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_132___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_132___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_133___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_133___stage___block_6_inside;
reg  [0:0] _d___pip_5160_1_134___stage___block_6_inside;
reg  [0:0] _q___pip_5160_1_134___stage___block_6_inside;
reg signed [23:0] _d___pip_5160_1_0___stage___block_6_view_x;
reg signed [23:0] _q___pip_5160_1_0___stage___block_6_view_x;
reg signed [23:0] _d___pip_5160_1_1___stage___block_6_view_x;
reg signed [23:0] _q___pip_5160_1_1___stage___block_6_view_x;
reg signed [23:0] _d___pip_5160_1_2___stage___block_6_view_x;
reg signed [23:0] _q___pip_5160_1_2___stage___block_6_view_x;
reg signed [23:0] _d___pip_5160_1_3___stage___block_6_view_x;
reg signed [23:0] _q___pip_5160_1_3___stage___block_6_view_x;
reg signed [23:0] _d___pip_5160_1_0___stage___block_6_view_y;
reg signed [23:0] _q___pip_5160_1_0___stage___block_6_view_y;
reg signed [23:0] _d___pip_5160_1_1___stage___block_6_view_y;
reg signed [23:0] _q___pip_5160_1_1___stage___block_6_view_y;
reg signed [23:0] _d___pip_5160_1_2___stage___block_6_view_y;
reg signed [23:0] _q___pip_5160_1_2___stage___block_6_view_y;
reg signed [23:0] _d___pip_5160_1_3___stage___block_6_view_y;
reg signed [23:0] _q___pip_5160_1_3___stage___block_6_view_y;
reg signed [23:0] _d___pip_5160_1_4___stage___block_6_view_y;
reg signed [23:0] _q___pip_5160_1_4___stage___block_6_view_y;
reg signed [23:0] _d___pip_5160_1_0___stage___block_6_view_z;
reg signed [23:0] _q___pip_5160_1_0___stage___block_6_view_z;
reg signed [23:0] _d___pip_5160_1_1___stage___block_6_view_z;
reg signed [23:0] _q___pip_5160_1_1___stage___block_6_view_z;
reg signed [23:0] _d___pip_5160_1_2___stage___block_6_view_z;
reg signed [23:0] _q___pip_5160_1_2___stage___block_6_view_z;
reg signed [23:0] _d___pip_5160_1_3___stage___block_6_view_z;
reg signed [23:0] _q___pip_5160_1_3___stage___block_6_view_z;
reg  [13:0] _d___pip_5160_1_0___stage___block_6_vxsz;
reg  [13:0] _q___pip_5160_1_0___stage___block_6_vxsz;
reg  [13:0] _d___pip_5160_1_1___stage___block_6_vxsz;
reg  [13:0] _q___pip_5160_1_1___stage___block_6_vxsz;
reg  [13:0] _d___pip_5160_1_2___stage___block_6_vxsz;
reg  [13:0] _q___pip_5160_1_2___stage___block_6_vxsz;
reg  [13:0] _d___pip_5160_1_3___stage___block_6_vxsz;
reg  [13:0] _q___pip_5160_1_3___stage___block_6_vxsz;
reg  [13:0] _d___pip_5160_1_4___stage___block_6_vxsz;
reg  [13:0] _q___pip_5160_1_4___stage___block_6_vxsz;
reg  [13:0] _d___pip_5160_1_5___stage___block_6_vxsz;
reg  [13:0] _q___pip_5160_1_5___stage___block_6_vxsz;
reg  [13:0] _d___pip_5160_1_6___stage___block_6_vxsz;
reg  [13:0] _q___pip_5160_1_6___stage___block_6_vxsz;
reg signed [23:0] _d___pip_5160_1_1___stage___block_7_cs0;
reg signed [23:0] _q___pip_5160_1_1___stage___block_7_cs0;
reg signed [23:0] _d___pip_5160_1_2___stage___block_7_cs0;
reg signed [23:0] _q___pip_5160_1_2___stage___block_7_cs0;
reg signed [23:0] _d___pip_5160_1_3___stage___block_7_cs0;
reg signed [23:0] _q___pip_5160_1_3___stage___block_7_cs0;
reg signed [23:0] _d___pip_5160_1_1___stage___block_7_ss0;
reg signed [23:0] _q___pip_5160_1_1___stage___block_7_ss0;
reg signed [23:0] _d___pip_5160_1_2___stage___block_7_ss0;
reg signed [23:0] _q___pip_5160_1_2___stage___block_7_ss0;
reg signed [23:0] _d___pip_5160_1_3___stage___block_7_ss0;
reg signed [23:0] _q___pip_5160_1_3___stage___block_7_ss0;
reg  [7:0] _d_pix_r;
reg  [7:0] _q_pix_r;
reg  [7:0] _d_pix_g;
reg  [7:0] _q_pix_g;
reg  [7:0] _d_pix_b;
reg  [7:0] _q_pix_b;
reg  [1:0] _d__idx_fsm0,_q__idx_fsm0;
reg  _autorun = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_0,_q__idx_fsm___pip_5160_1_0;
wire _ready_fsm___pip_5160_1_0 = (_q__idx_fsm___pip_5160_1_0 == 1) || (_q__idx_fsm___pip_5160_1_0 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_0 = 0,_q__full_fsm___pip_5160_1_0 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_0 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_0 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_1,_q__idx_fsm___pip_5160_1_1;
wire _ready_fsm___pip_5160_1_1 = (_q__idx_fsm___pip_5160_1_1 == 1) || (_q__idx_fsm___pip_5160_1_1 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_1 = 0,_q__full_fsm___pip_5160_1_1 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_1 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_1 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_2,_q__idx_fsm___pip_5160_1_2;
wire _ready_fsm___pip_5160_1_2 = (_q__idx_fsm___pip_5160_1_2 == 1) || (_q__idx_fsm___pip_5160_1_2 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_2 = 0,_q__full_fsm___pip_5160_1_2 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_2 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_2 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_3,_q__idx_fsm___pip_5160_1_3;
wire _ready_fsm___pip_5160_1_3 = (_q__idx_fsm___pip_5160_1_3 == 1) || (_q__idx_fsm___pip_5160_1_3 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_3 = 0,_q__full_fsm___pip_5160_1_3 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_3 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_3 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_4,_q__idx_fsm___pip_5160_1_4;
wire _ready_fsm___pip_5160_1_4 = (_q__idx_fsm___pip_5160_1_4 == 1) || (_q__idx_fsm___pip_5160_1_4 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_4 = 0,_q__full_fsm___pip_5160_1_4 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_4 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_4 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_5,_q__idx_fsm___pip_5160_1_5;
wire _ready_fsm___pip_5160_1_5 = (_q__idx_fsm___pip_5160_1_5 == 1) || (_q__idx_fsm___pip_5160_1_5 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_5 = 0,_q__full_fsm___pip_5160_1_5 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_5 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_5 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_6,_q__idx_fsm___pip_5160_1_6;
wire _ready_fsm___pip_5160_1_6 = (_q__idx_fsm___pip_5160_1_6 == 1) || (_q__idx_fsm___pip_5160_1_6 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_6 = 0,_q__full_fsm___pip_5160_1_6 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_6 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_6 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_7,_q__idx_fsm___pip_5160_1_7;
wire _ready_fsm___pip_5160_1_7 = (_q__idx_fsm___pip_5160_1_7 == 1) || (_q__idx_fsm___pip_5160_1_7 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_7 = 0,_q__full_fsm___pip_5160_1_7 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_7 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_7 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_8,_q__idx_fsm___pip_5160_1_8;
wire _ready_fsm___pip_5160_1_8 = (_q__idx_fsm___pip_5160_1_8 == 1) || (_q__idx_fsm___pip_5160_1_8 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_8 = 0,_q__full_fsm___pip_5160_1_8 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_8 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_8 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_9,_q__idx_fsm___pip_5160_1_9;
wire _ready_fsm___pip_5160_1_9 = (_q__idx_fsm___pip_5160_1_9 == 1) || (_q__idx_fsm___pip_5160_1_9 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_9 = 0,_q__full_fsm___pip_5160_1_9 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_9 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_9 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_10,_q__idx_fsm___pip_5160_1_10;
wire _ready_fsm___pip_5160_1_10 = (_q__idx_fsm___pip_5160_1_10 == 1) || (_q__idx_fsm___pip_5160_1_10 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_10 = 0,_q__full_fsm___pip_5160_1_10 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_10 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_10 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_11,_q__idx_fsm___pip_5160_1_11;
wire _ready_fsm___pip_5160_1_11 = (_q__idx_fsm___pip_5160_1_11 == 1) || (_q__idx_fsm___pip_5160_1_11 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_11 = 0,_q__full_fsm___pip_5160_1_11 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_11 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_11 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_12,_q__idx_fsm___pip_5160_1_12;
wire _ready_fsm___pip_5160_1_12 = (_q__idx_fsm___pip_5160_1_12 == 1) || (_q__idx_fsm___pip_5160_1_12 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_12 = 0,_q__full_fsm___pip_5160_1_12 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_12 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_12 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_13,_q__idx_fsm___pip_5160_1_13;
wire _ready_fsm___pip_5160_1_13 = (_q__idx_fsm___pip_5160_1_13 == 1) || (_q__idx_fsm___pip_5160_1_13 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_13 = 0,_q__full_fsm___pip_5160_1_13 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_13 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_13 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_14,_q__idx_fsm___pip_5160_1_14;
wire _ready_fsm___pip_5160_1_14 = (_q__idx_fsm___pip_5160_1_14 == 1) || (_q__idx_fsm___pip_5160_1_14 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_14 = 0,_q__full_fsm___pip_5160_1_14 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_14 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_14 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_15,_q__idx_fsm___pip_5160_1_15;
wire _ready_fsm___pip_5160_1_15 = (_q__idx_fsm___pip_5160_1_15 == 1) || (_q__idx_fsm___pip_5160_1_15 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_15 = 0,_q__full_fsm___pip_5160_1_15 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_15 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_15 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_16,_q__idx_fsm___pip_5160_1_16;
wire _ready_fsm___pip_5160_1_16 = (_q__idx_fsm___pip_5160_1_16 == 1) || (_q__idx_fsm___pip_5160_1_16 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_16 = 0,_q__full_fsm___pip_5160_1_16 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_16 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_16 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_17,_q__idx_fsm___pip_5160_1_17;
wire _ready_fsm___pip_5160_1_17 = (_q__idx_fsm___pip_5160_1_17 == 1) || (_q__idx_fsm___pip_5160_1_17 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_17 = 0,_q__full_fsm___pip_5160_1_17 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_17 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_17 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_18,_q__idx_fsm___pip_5160_1_18;
wire _ready_fsm___pip_5160_1_18 = (_q__idx_fsm___pip_5160_1_18 == 1) || (_q__idx_fsm___pip_5160_1_18 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_18 = 0,_q__full_fsm___pip_5160_1_18 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_18 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_18 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_19,_q__idx_fsm___pip_5160_1_19;
wire _ready_fsm___pip_5160_1_19 = (_q__idx_fsm___pip_5160_1_19 == 1) || (_q__idx_fsm___pip_5160_1_19 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_19 = 0,_q__full_fsm___pip_5160_1_19 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_19 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_19 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_20,_q__idx_fsm___pip_5160_1_20;
wire _ready_fsm___pip_5160_1_20 = (_q__idx_fsm___pip_5160_1_20 == 1) || (_q__idx_fsm___pip_5160_1_20 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_20 = 0,_q__full_fsm___pip_5160_1_20 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_20 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_20 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_21,_q__idx_fsm___pip_5160_1_21;
wire _ready_fsm___pip_5160_1_21 = (_q__idx_fsm___pip_5160_1_21 == 1) || (_q__idx_fsm___pip_5160_1_21 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_21 = 0,_q__full_fsm___pip_5160_1_21 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_21 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_21 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_22,_q__idx_fsm___pip_5160_1_22;
wire _ready_fsm___pip_5160_1_22 = (_q__idx_fsm___pip_5160_1_22 == 1) || (_q__idx_fsm___pip_5160_1_22 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_22 = 0,_q__full_fsm___pip_5160_1_22 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_22 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_22 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_23,_q__idx_fsm___pip_5160_1_23;
wire _ready_fsm___pip_5160_1_23 = (_q__idx_fsm___pip_5160_1_23 == 1) || (_q__idx_fsm___pip_5160_1_23 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_23 = 0,_q__full_fsm___pip_5160_1_23 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_23 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_23 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_24,_q__idx_fsm___pip_5160_1_24;
wire _ready_fsm___pip_5160_1_24 = (_q__idx_fsm___pip_5160_1_24 == 1) || (_q__idx_fsm___pip_5160_1_24 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_24 = 0,_q__full_fsm___pip_5160_1_24 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_24 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_24 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_25,_q__idx_fsm___pip_5160_1_25;
wire _ready_fsm___pip_5160_1_25 = (_q__idx_fsm___pip_5160_1_25 == 1) || (_q__idx_fsm___pip_5160_1_25 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_25 = 0,_q__full_fsm___pip_5160_1_25 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_25 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_25 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_26,_q__idx_fsm___pip_5160_1_26;
wire _ready_fsm___pip_5160_1_26 = (_q__idx_fsm___pip_5160_1_26 == 1) || (_q__idx_fsm___pip_5160_1_26 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_26 = 0,_q__full_fsm___pip_5160_1_26 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_26 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_26 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_27,_q__idx_fsm___pip_5160_1_27;
wire _ready_fsm___pip_5160_1_27 = (_q__idx_fsm___pip_5160_1_27 == 1) || (_q__idx_fsm___pip_5160_1_27 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_27 = 0,_q__full_fsm___pip_5160_1_27 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_27 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_27 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_28,_q__idx_fsm___pip_5160_1_28;
wire _ready_fsm___pip_5160_1_28 = (_q__idx_fsm___pip_5160_1_28 == 1) || (_q__idx_fsm___pip_5160_1_28 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_28 = 0,_q__full_fsm___pip_5160_1_28 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_28 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_28 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_29,_q__idx_fsm___pip_5160_1_29;
wire _ready_fsm___pip_5160_1_29 = (_q__idx_fsm___pip_5160_1_29 == 1) || (_q__idx_fsm___pip_5160_1_29 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_29 = 0,_q__full_fsm___pip_5160_1_29 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_29 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_29 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_30,_q__idx_fsm___pip_5160_1_30;
wire _ready_fsm___pip_5160_1_30 = (_q__idx_fsm___pip_5160_1_30 == 1) || (_q__idx_fsm___pip_5160_1_30 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_30 = 0,_q__full_fsm___pip_5160_1_30 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_30 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_30 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_31,_q__idx_fsm___pip_5160_1_31;
wire _ready_fsm___pip_5160_1_31 = (_q__idx_fsm___pip_5160_1_31 == 1) || (_q__idx_fsm___pip_5160_1_31 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_31 = 0,_q__full_fsm___pip_5160_1_31 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_31 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_31 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_32,_q__idx_fsm___pip_5160_1_32;
wire _ready_fsm___pip_5160_1_32 = (_q__idx_fsm___pip_5160_1_32 == 1) || (_q__idx_fsm___pip_5160_1_32 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_32 = 0,_q__full_fsm___pip_5160_1_32 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_32 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_32 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_33,_q__idx_fsm___pip_5160_1_33;
wire _ready_fsm___pip_5160_1_33 = (_q__idx_fsm___pip_5160_1_33 == 1) || (_q__idx_fsm___pip_5160_1_33 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_33 = 0,_q__full_fsm___pip_5160_1_33 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_33 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_33 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_34,_q__idx_fsm___pip_5160_1_34;
wire _ready_fsm___pip_5160_1_34 = (_q__idx_fsm___pip_5160_1_34 == 1) || (_q__idx_fsm___pip_5160_1_34 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_34 = 0,_q__full_fsm___pip_5160_1_34 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_34 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_34 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_35,_q__idx_fsm___pip_5160_1_35;
wire _ready_fsm___pip_5160_1_35 = (_q__idx_fsm___pip_5160_1_35 == 1) || (_q__idx_fsm___pip_5160_1_35 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_35 = 0,_q__full_fsm___pip_5160_1_35 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_35 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_35 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_36,_q__idx_fsm___pip_5160_1_36;
wire _ready_fsm___pip_5160_1_36 = (_q__idx_fsm___pip_5160_1_36 == 1) || (_q__idx_fsm___pip_5160_1_36 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_36 = 0,_q__full_fsm___pip_5160_1_36 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_36 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_36 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_37,_q__idx_fsm___pip_5160_1_37;
wire _ready_fsm___pip_5160_1_37 = (_q__idx_fsm___pip_5160_1_37 == 1) || (_q__idx_fsm___pip_5160_1_37 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_37 = 0,_q__full_fsm___pip_5160_1_37 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_37 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_37 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_38,_q__idx_fsm___pip_5160_1_38;
wire _ready_fsm___pip_5160_1_38 = (_q__idx_fsm___pip_5160_1_38 == 1) || (_q__idx_fsm___pip_5160_1_38 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_38 = 0,_q__full_fsm___pip_5160_1_38 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_38 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_38 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_39,_q__idx_fsm___pip_5160_1_39;
wire _ready_fsm___pip_5160_1_39 = (_q__idx_fsm___pip_5160_1_39 == 1) || (_q__idx_fsm___pip_5160_1_39 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_39 = 0,_q__full_fsm___pip_5160_1_39 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_39 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_39 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_40,_q__idx_fsm___pip_5160_1_40;
wire _ready_fsm___pip_5160_1_40 = (_q__idx_fsm___pip_5160_1_40 == 1) || (_q__idx_fsm___pip_5160_1_40 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_40 = 0,_q__full_fsm___pip_5160_1_40 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_40 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_40 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_41,_q__idx_fsm___pip_5160_1_41;
wire _ready_fsm___pip_5160_1_41 = (_q__idx_fsm___pip_5160_1_41 == 1) || (_q__idx_fsm___pip_5160_1_41 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_41 = 0,_q__full_fsm___pip_5160_1_41 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_41 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_41 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_42,_q__idx_fsm___pip_5160_1_42;
wire _ready_fsm___pip_5160_1_42 = (_q__idx_fsm___pip_5160_1_42 == 1) || (_q__idx_fsm___pip_5160_1_42 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_42 = 0,_q__full_fsm___pip_5160_1_42 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_42 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_42 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_43,_q__idx_fsm___pip_5160_1_43;
wire _ready_fsm___pip_5160_1_43 = (_q__idx_fsm___pip_5160_1_43 == 1) || (_q__idx_fsm___pip_5160_1_43 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_43 = 0,_q__full_fsm___pip_5160_1_43 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_43 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_43 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_44,_q__idx_fsm___pip_5160_1_44;
wire _ready_fsm___pip_5160_1_44 = (_q__idx_fsm___pip_5160_1_44 == 1) || (_q__idx_fsm___pip_5160_1_44 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_44 = 0,_q__full_fsm___pip_5160_1_44 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_44 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_44 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_45,_q__idx_fsm___pip_5160_1_45;
wire _ready_fsm___pip_5160_1_45 = (_q__idx_fsm___pip_5160_1_45 == 1) || (_q__idx_fsm___pip_5160_1_45 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_45 = 0,_q__full_fsm___pip_5160_1_45 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_45 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_45 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_46,_q__idx_fsm___pip_5160_1_46;
wire _ready_fsm___pip_5160_1_46 = (_q__idx_fsm___pip_5160_1_46 == 1) || (_q__idx_fsm___pip_5160_1_46 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_46 = 0,_q__full_fsm___pip_5160_1_46 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_46 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_46 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_47,_q__idx_fsm___pip_5160_1_47;
wire _ready_fsm___pip_5160_1_47 = (_q__idx_fsm___pip_5160_1_47 == 1) || (_q__idx_fsm___pip_5160_1_47 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_47 = 0,_q__full_fsm___pip_5160_1_47 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_47 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_47 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_48,_q__idx_fsm___pip_5160_1_48;
wire _ready_fsm___pip_5160_1_48 = (_q__idx_fsm___pip_5160_1_48 == 1) || (_q__idx_fsm___pip_5160_1_48 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_48 = 0,_q__full_fsm___pip_5160_1_48 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_48 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_48 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_49,_q__idx_fsm___pip_5160_1_49;
wire _ready_fsm___pip_5160_1_49 = (_q__idx_fsm___pip_5160_1_49 == 1) || (_q__idx_fsm___pip_5160_1_49 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_49 = 0,_q__full_fsm___pip_5160_1_49 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_49 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_49 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_50,_q__idx_fsm___pip_5160_1_50;
wire _ready_fsm___pip_5160_1_50 = (_q__idx_fsm___pip_5160_1_50 == 1) || (_q__idx_fsm___pip_5160_1_50 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_50 = 0,_q__full_fsm___pip_5160_1_50 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_50 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_50 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_51,_q__idx_fsm___pip_5160_1_51;
wire _ready_fsm___pip_5160_1_51 = (_q__idx_fsm___pip_5160_1_51 == 1) || (_q__idx_fsm___pip_5160_1_51 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_51 = 0,_q__full_fsm___pip_5160_1_51 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_51 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_51 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_52,_q__idx_fsm___pip_5160_1_52;
wire _ready_fsm___pip_5160_1_52 = (_q__idx_fsm___pip_5160_1_52 == 1) || (_q__idx_fsm___pip_5160_1_52 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_52 = 0,_q__full_fsm___pip_5160_1_52 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_52 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_52 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_53,_q__idx_fsm___pip_5160_1_53;
wire _ready_fsm___pip_5160_1_53 = (_q__idx_fsm___pip_5160_1_53 == 1) || (_q__idx_fsm___pip_5160_1_53 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_53 = 0,_q__full_fsm___pip_5160_1_53 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_53 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_53 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_54,_q__idx_fsm___pip_5160_1_54;
wire _ready_fsm___pip_5160_1_54 = (_q__idx_fsm___pip_5160_1_54 == 1) || (_q__idx_fsm___pip_5160_1_54 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_54 = 0,_q__full_fsm___pip_5160_1_54 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_54 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_54 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_55,_q__idx_fsm___pip_5160_1_55;
wire _ready_fsm___pip_5160_1_55 = (_q__idx_fsm___pip_5160_1_55 == 1) || (_q__idx_fsm___pip_5160_1_55 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_55 = 0,_q__full_fsm___pip_5160_1_55 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_55 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_55 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_56,_q__idx_fsm___pip_5160_1_56;
wire _ready_fsm___pip_5160_1_56 = (_q__idx_fsm___pip_5160_1_56 == 1) || (_q__idx_fsm___pip_5160_1_56 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_56 = 0,_q__full_fsm___pip_5160_1_56 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_56 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_56 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_57,_q__idx_fsm___pip_5160_1_57;
wire _ready_fsm___pip_5160_1_57 = (_q__idx_fsm___pip_5160_1_57 == 1) || (_q__idx_fsm___pip_5160_1_57 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_57 = 0,_q__full_fsm___pip_5160_1_57 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_57 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_57 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_58,_q__idx_fsm___pip_5160_1_58;
wire _ready_fsm___pip_5160_1_58 = (_q__idx_fsm___pip_5160_1_58 == 1) || (_q__idx_fsm___pip_5160_1_58 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_58 = 0,_q__full_fsm___pip_5160_1_58 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_58 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_58 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_59,_q__idx_fsm___pip_5160_1_59;
wire _ready_fsm___pip_5160_1_59 = (_q__idx_fsm___pip_5160_1_59 == 1) || (_q__idx_fsm___pip_5160_1_59 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_59 = 0,_q__full_fsm___pip_5160_1_59 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_59 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_59 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_60,_q__idx_fsm___pip_5160_1_60;
wire _ready_fsm___pip_5160_1_60 = (_q__idx_fsm___pip_5160_1_60 == 1) || (_q__idx_fsm___pip_5160_1_60 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_60 = 0,_q__full_fsm___pip_5160_1_60 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_60 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_60 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_61,_q__idx_fsm___pip_5160_1_61;
wire _ready_fsm___pip_5160_1_61 = (_q__idx_fsm___pip_5160_1_61 == 1) || (_q__idx_fsm___pip_5160_1_61 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_61 = 0,_q__full_fsm___pip_5160_1_61 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_61 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_61 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_62,_q__idx_fsm___pip_5160_1_62;
wire _ready_fsm___pip_5160_1_62 = (_q__idx_fsm___pip_5160_1_62 == 1) || (_q__idx_fsm___pip_5160_1_62 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_62 = 0,_q__full_fsm___pip_5160_1_62 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_62 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_62 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_63,_q__idx_fsm___pip_5160_1_63;
wire _ready_fsm___pip_5160_1_63 = (_q__idx_fsm___pip_5160_1_63 == 1) || (_q__idx_fsm___pip_5160_1_63 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_63 = 0,_q__full_fsm___pip_5160_1_63 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_63 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_63 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_64,_q__idx_fsm___pip_5160_1_64;
wire _ready_fsm___pip_5160_1_64 = (_q__idx_fsm___pip_5160_1_64 == 1) || (_q__idx_fsm___pip_5160_1_64 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_64 = 0,_q__full_fsm___pip_5160_1_64 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_64 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_64 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_65,_q__idx_fsm___pip_5160_1_65;
wire _ready_fsm___pip_5160_1_65 = (_q__idx_fsm___pip_5160_1_65 == 1) || (_q__idx_fsm___pip_5160_1_65 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_65 = 0,_q__full_fsm___pip_5160_1_65 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_65 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_65 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_66,_q__idx_fsm___pip_5160_1_66;
wire _ready_fsm___pip_5160_1_66 = (_q__idx_fsm___pip_5160_1_66 == 1) || (_q__idx_fsm___pip_5160_1_66 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_66 = 0,_q__full_fsm___pip_5160_1_66 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_66 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_66 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_67,_q__idx_fsm___pip_5160_1_67;
wire _ready_fsm___pip_5160_1_67 = (_q__idx_fsm___pip_5160_1_67 == 1) || (_q__idx_fsm___pip_5160_1_67 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_67 = 0,_q__full_fsm___pip_5160_1_67 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_67 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_67 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_68,_q__idx_fsm___pip_5160_1_68;
wire _ready_fsm___pip_5160_1_68 = (_q__idx_fsm___pip_5160_1_68 == 1) || (_q__idx_fsm___pip_5160_1_68 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_68 = 0,_q__full_fsm___pip_5160_1_68 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_68 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_68 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_69,_q__idx_fsm___pip_5160_1_69;
wire _ready_fsm___pip_5160_1_69 = (_q__idx_fsm___pip_5160_1_69 == 1) || (_q__idx_fsm___pip_5160_1_69 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_69 = 0,_q__full_fsm___pip_5160_1_69 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_69 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_69 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_70,_q__idx_fsm___pip_5160_1_70;
wire _ready_fsm___pip_5160_1_70 = (_q__idx_fsm___pip_5160_1_70 == 1) || (_q__idx_fsm___pip_5160_1_70 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_70 = 0,_q__full_fsm___pip_5160_1_70 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_70 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_70 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_71,_q__idx_fsm___pip_5160_1_71;
wire _ready_fsm___pip_5160_1_71 = (_q__idx_fsm___pip_5160_1_71 == 1) || (_q__idx_fsm___pip_5160_1_71 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_71 = 0,_q__full_fsm___pip_5160_1_71 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_71 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_71 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_72,_q__idx_fsm___pip_5160_1_72;
wire _ready_fsm___pip_5160_1_72 = (_q__idx_fsm___pip_5160_1_72 == 1) || (_q__idx_fsm___pip_5160_1_72 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_72 = 0,_q__full_fsm___pip_5160_1_72 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_72 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_72 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_73,_q__idx_fsm___pip_5160_1_73;
wire _ready_fsm___pip_5160_1_73 = (_q__idx_fsm___pip_5160_1_73 == 1) || (_q__idx_fsm___pip_5160_1_73 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_73 = 0,_q__full_fsm___pip_5160_1_73 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_73 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_73 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_74,_q__idx_fsm___pip_5160_1_74;
wire _ready_fsm___pip_5160_1_74 = (_q__idx_fsm___pip_5160_1_74 == 1) || (_q__idx_fsm___pip_5160_1_74 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_74 = 0,_q__full_fsm___pip_5160_1_74 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_74 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_74 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_75,_q__idx_fsm___pip_5160_1_75;
wire _ready_fsm___pip_5160_1_75 = (_q__idx_fsm___pip_5160_1_75 == 1) || (_q__idx_fsm___pip_5160_1_75 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_75 = 0,_q__full_fsm___pip_5160_1_75 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_75 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_75 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_76,_q__idx_fsm___pip_5160_1_76;
wire _ready_fsm___pip_5160_1_76 = (_q__idx_fsm___pip_5160_1_76 == 1) || (_q__idx_fsm___pip_5160_1_76 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_76 = 0,_q__full_fsm___pip_5160_1_76 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_76 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_76 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_77,_q__idx_fsm___pip_5160_1_77;
wire _ready_fsm___pip_5160_1_77 = (_q__idx_fsm___pip_5160_1_77 == 1) || (_q__idx_fsm___pip_5160_1_77 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_77 = 0,_q__full_fsm___pip_5160_1_77 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_77 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_77 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_78,_q__idx_fsm___pip_5160_1_78;
wire _ready_fsm___pip_5160_1_78 = (_q__idx_fsm___pip_5160_1_78 == 1) || (_q__idx_fsm___pip_5160_1_78 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_78 = 0,_q__full_fsm___pip_5160_1_78 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_78 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_78 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_79,_q__idx_fsm___pip_5160_1_79;
wire _ready_fsm___pip_5160_1_79 = (_q__idx_fsm___pip_5160_1_79 == 1) || (_q__idx_fsm___pip_5160_1_79 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_79 = 0,_q__full_fsm___pip_5160_1_79 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_79 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_79 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_80,_q__idx_fsm___pip_5160_1_80;
wire _ready_fsm___pip_5160_1_80 = (_q__idx_fsm___pip_5160_1_80 == 1) || (_q__idx_fsm___pip_5160_1_80 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_80 = 0,_q__full_fsm___pip_5160_1_80 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_80 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_80 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_81,_q__idx_fsm___pip_5160_1_81;
wire _ready_fsm___pip_5160_1_81 = (_q__idx_fsm___pip_5160_1_81 == 1) || (_q__idx_fsm___pip_5160_1_81 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_81 = 0,_q__full_fsm___pip_5160_1_81 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_81 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_81 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_82,_q__idx_fsm___pip_5160_1_82;
wire _ready_fsm___pip_5160_1_82 = (_q__idx_fsm___pip_5160_1_82 == 1) || (_q__idx_fsm___pip_5160_1_82 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_82 = 0,_q__full_fsm___pip_5160_1_82 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_82 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_82 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_83,_q__idx_fsm___pip_5160_1_83;
wire _ready_fsm___pip_5160_1_83 = (_q__idx_fsm___pip_5160_1_83 == 1) || (_q__idx_fsm___pip_5160_1_83 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_83 = 0,_q__full_fsm___pip_5160_1_83 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_83 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_83 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_84,_q__idx_fsm___pip_5160_1_84;
wire _ready_fsm___pip_5160_1_84 = (_q__idx_fsm___pip_5160_1_84 == 1) || (_q__idx_fsm___pip_5160_1_84 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_84 = 0,_q__full_fsm___pip_5160_1_84 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_84 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_84 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_85,_q__idx_fsm___pip_5160_1_85;
wire _ready_fsm___pip_5160_1_85 = (_q__idx_fsm___pip_5160_1_85 == 1) || (_q__idx_fsm___pip_5160_1_85 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_85 = 0,_q__full_fsm___pip_5160_1_85 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_85 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_85 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_86,_q__idx_fsm___pip_5160_1_86;
wire _ready_fsm___pip_5160_1_86 = (_q__idx_fsm___pip_5160_1_86 == 1) || (_q__idx_fsm___pip_5160_1_86 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_86 = 0,_q__full_fsm___pip_5160_1_86 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_86 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_86 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_87,_q__idx_fsm___pip_5160_1_87;
wire _ready_fsm___pip_5160_1_87 = (_q__idx_fsm___pip_5160_1_87 == 1) || (_q__idx_fsm___pip_5160_1_87 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_87 = 0,_q__full_fsm___pip_5160_1_87 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_87 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_87 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_88,_q__idx_fsm___pip_5160_1_88;
wire _ready_fsm___pip_5160_1_88 = (_q__idx_fsm___pip_5160_1_88 == 1) || (_q__idx_fsm___pip_5160_1_88 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_88 = 0,_q__full_fsm___pip_5160_1_88 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_88 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_88 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_89,_q__idx_fsm___pip_5160_1_89;
wire _ready_fsm___pip_5160_1_89 = (_q__idx_fsm___pip_5160_1_89 == 1) || (_q__idx_fsm___pip_5160_1_89 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_89 = 0,_q__full_fsm___pip_5160_1_89 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_89 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_89 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_90,_q__idx_fsm___pip_5160_1_90;
wire _ready_fsm___pip_5160_1_90 = (_q__idx_fsm___pip_5160_1_90 == 1) || (_q__idx_fsm___pip_5160_1_90 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_90 = 0,_q__full_fsm___pip_5160_1_90 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_90 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_90 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_91,_q__idx_fsm___pip_5160_1_91;
wire _ready_fsm___pip_5160_1_91 = (_q__idx_fsm___pip_5160_1_91 == 1) || (_q__idx_fsm___pip_5160_1_91 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_91 = 0,_q__full_fsm___pip_5160_1_91 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_91 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_91 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_92,_q__idx_fsm___pip_5160_1_92;
wire _ready_fsm___pip_5160_1_92 = (_q__idx_fsm___pip_5160_1_92 == 1) || (_q__idx_fsm___pip_5160_1_92 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_92 = 0,_q__full_fsm___pip_5160_1_92 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_92 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_92 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_93,_q__idx_fsm___pip_5160_1_93;
wire _ready_fsm___pip_5160_1_93 = (_q__idx_fsm___pip_5160_1_93 == 1) || (_q__idx_fsm___pip_5160_1_93 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_93 = 0,_q__full_fsm___pip_5160_1_93 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_93 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_93 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_94,_q__idx_fsm___pip_5160_1_94;
wire _ready_fsm___pip_5160_1_94 = (_q__idx_fsm___pip_5160_1_94 == 1) || (_q__idx_fsm___pip_5160_1_94 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_94 = 0,_q__full_fsm___pip_5160_1_94 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_94 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_94 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_95,_q__idx_fsm___pip_5160_1_95;
wire _ready_fsm___pip_5160_1_95 = (_q__idx_fsm___pip_5160_1_95 == 1) || (_q__idx_fsm___pip_5160_1_95 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_95 = 0,_q__full_fsm___pip_5160_1_95 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_95 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_95 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_96,_q__idx_fsm___pip_5160_1_96;
wire _ready_fsm___pip_5160_1_96 = (_q__idx_fsm___pip_5160_1_96 == 1) || (_q__idx_fsm___pip_5160_1_96 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_96 = 0,_q__full_fsm___pip_5160_1_96 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_96 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_96 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_97,_q__idx_fsm___pip_5160_1_97;
wire _ready_fsm___pip_5160_1_97 = (_q__idx_fsm___pip_5160_1_97 == 1) || (_q__idx_fsm___pip_5160_1_97 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_97 = 0,_q__full_fsm___pip_5160_1_97 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_97 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_97 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_98,_q__idx_fsm___pip_5160_1_98;
wire _ready_fsm___pip_5160_1_98 = (_q__idx_fsm___pip_5160_1_98 == 1) || (_q__idx_fsm___pip_5160_1_98 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_98 = 0,_q__full_fsm___pip_5160_1_98 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_98 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_98 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_99,_q__idx_fsm___pip_5160_1_99;
wire _ready_fsm___pip_5160_1_99 = (_q__idx_fsm___pip_5160_1_99 == 1) || (_q__idx_fsm___pip_5160_1_99 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_99 = 0,_q__full_fsm___pip_5160_1_99 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_99 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_99 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_100,_q__idx_fsm___pip_5160_1_100;
wire _ready_fsm___pip_5160_1_100 = (_q__idx_fsm___pip_5160_1_100 == 1) || (_q__idx_fsm___pip_5160_1_100 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_100 = 0,_q__full_fsm___pip_5160_1_100 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_100 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_100 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_101,_q__idx_fsm___pip_5160_1_101;
wire _ready_fsm___pip_5160_1_101 = (_q__idx_fsm___pip_5160_1_101 == 1) || (_q__idx_fsm___pip_5160_1_101 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_101 = 0,_q__full_fsm___pip_5160_1_101 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_101 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_101 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_102,_q__idx_fsm___pip_5160_1_102;
wire _ready_fsm___pip_5160_1_102 = (_q__idx_fsm___pip_5160_1_102 == 1) || (_q__idx_fsm___pip_5160_1_102 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_102 = 0,_q__full_fsm___pip_5160_1_102 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_102 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_102 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_103,_q__idx_fsm___pip_5160_1_103;
wire _ready_fsm___pip_5160_1_103 = (_q__idx_fsm___pip_5160_1_103 == 1) || (_q__idx_fsm___pip_5160_1_103 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_103 = 0,_q__full_fsm___pip_5160_1_103 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_103 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_103 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_104,_q__idx_fsm___pip_5160_1_104;
wire _ready_fsm___pip_5160_1_104 = (_q__idx_fsm___pip_5160_1_104 == 1) || (_q__idx_fsm___pip_5160_1_104 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_104 = 0,_q__full_fsm___pip_5160_1_104 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_104 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_104 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_105,_q__idx_fsm___pip_5160_1_105;
wire _ready_fsm___pip_5160_1_105 = (_q__idx_fsm___pip_5160_1_105 == 1) || (_q__idx_fsm___pip_5160_1_105 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_105 = 0,_q__full_fsm___pip_5160_1_105 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_105 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_105 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_106,_q__idx_fsm___pip_5160_1_106;
wire _ready_fsm___pip_5160_1_106 = (_q__idx_fsm___pip_5160_1_106 == 1) || (_q__idx_fsm___pip_5160_1_106 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_106 = 0,_q__full_fsm___pip_5160_1_106 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_106 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_106 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_107,_q__idx_fsm___pip_5160_1_107;
wire _ready_fsm___pip_5160_1_107 = (_q__idx_fsm___pip_5160_1_107 == 1) || (_q__idx_fsm___pip_5160_1_107 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_107 = 0,_q__full_fsm___pip_5160_1_107 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_107 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_107 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_108,_q__idx_fsm___pip_5160_1_108;
wire _ready_fsm___pip_5160_1_108 = (_q__idx_fsm___pip_5160_1_108 == 1) || (_q__idx_fsm___pip_5160_1_108 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_108 = 0,_q__full_fsm___pip_5160_1_108 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_108 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_108 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_109,_q__idx_fsm___pip_5160_1_109;
wire _ready_fsm___pip_5160_1_109 = (_q__idx_fsm___pip_5160_1_109 == 1) || (_q__idx_fsm___pip_5160_1_109 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_109 = 0,_q__full_fsm___pip_5160_1_109 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_109 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_109 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_110,_q__idx_fsm___pip_5160_1_110;
wire _ready_fsm___pip_5160_1_110 = (_q__idx_fsm___pip_5160_1_110 == 1) || (_q__idx_fsm___pip_5160_1_110 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_110 = 0,_q__full_fsm___pip_5160_1_110 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_110 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_110 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_111,_q__idx_fsm___pip_5160_1_111;
wire _ready_fsm___pip_5160_1_111 = (_q__idx_fsm___pip_5160_1_111 == 1) || (_q__idx_fsm___pip_5160_1_111 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_111 = 0,_q__full_fsm___pip_5160_1_111 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_111 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_111 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_112,_q__idx_fsm___pip_5160_1_112;
wire _ready_fsm___pip_5160_1_112 = (_q__idx_fsm___pip_5160_1_112 == 1) || (_q__idx_fsm___pip_5160_1_112 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_112 = 0,_q__full_fsm___pip_5160_1_112 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_112 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_112 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_113,_q__idx_fsm___pip_5160_1_113;
wire _ready_fsm___pip_5160_1_113 = (_q__idx_fsm___pip_5160_1_113 == 1) || (_q__idx_fsm___pip_5160_1_113 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_113 = 0,_q__full_fsm___pip_5160_1_113 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_113 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_113 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_114,_q__idx_fsm___pip_5160_1_114;
wire _ready_fsm___pip_5160_1_114 = (_q__idx_fsm___pip_5160_1_114 == 1) || (_q__idx_fsm___pip_5160_1_114 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_114 = 0,_q__full_fsm___pip_5160_1_114 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_114 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_114 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_115,_q__idx_fsm___pip_5160_1_115;
wire _ready_fsm___pip_5160_1_115 = (_q__idx_fsm___pip_5160_1_115 == 1) || (_q__idx_fsm___pip_5160_1_115 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_115 = 0,_q__full_fsm___pip_5160_1_115 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_115 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_115 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_116,_q__idx_fsm___pip_5160_1_116;
wire _ready_fsm___pip_5160_1_116 = (_q__idx_fsm___pip_5160_1_116 == 1) || (_q__idx_fsm___pip_5160_1_116 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_116 = 0,_q__full_fsm___pip_5160_1_116 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_116 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_116 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_117,_q__idx_fsm___pip_5160_1_117;
wire _ready_fsm___pip_5160_1_117 = (_q__idx_fsm___pip_5160_1_117 == 1) || (_q__idx_fsm___pip_5160_1_117 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_117 = 0,_q__full_fsm___pip_5160_1_117 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_117 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_117 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_118,_q__idx_fsm___pip_5160_1_118;
wire _ready_fsm___pip_5160_1_118 = (_q__idx_fsm___pip_5160_1_118 == 1) || (_q__idx_fsm___pip_5160_1_118 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_118 = 0,_q__full_fsm___pip_5160_1_118 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_118 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_118 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_119,_q__idx_fsm___pip_5160_1_119;
wire _ready_fsm___pip_5160_1_119 = (_q__idx_fsm___pip_5160_1_119 == 1) || (_q__idx_fsm___pip_5160_1_119 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_119 = 0,_q__full_fsm___pip_5160_1_119 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_119 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_119 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_120,_q__idx_fsm___pip_5160_1_120;
wire _ready_fsm___pip_5160_1_120 = (_q__idx_fsm___pip_5160_1_120 == 1) || (_q__idx_fsm___pip_5160_1_120 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_120 = 0,_q__full_fsm___pip_5160_1_120 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_120 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_120 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_121,_q__idx_fsm___pip_5160_1_121;
wire _ready_fsm___pip_5160_1_121 = (_q__idx_fsm___pip_5160_1_121 == 1) || (_q__idx_fsm___pip_5160_1_121 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_121 = 0,_q__full_fsm___pip_5160_1_121 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_121 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_121 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_122,_q__idx_fsm___pip_5160_1_122;
wire _ready_fsm___pip_5160_1_122 = (_q__idx_fsm___pip_5160_1_122 == 1) || (_q__idx_fsm___pip_5160_1_122 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_122 = 0,_q__full_fsm___pip_5160_1_122 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_122 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_122 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_123,_q__idx_fsm___pip_5160_1_123;
wire _ready_fsm___pip_5160_1_123 = (_q__idx_fsm___pip_5160_1_123 == 1) || (_q__idx_fsm___pip_5160_1_123 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_123 = 0,_q__full_fsm___pip_5160_1_123 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_123 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_123 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_124,_q__idx_fsm___pip_5160_1_124;
wire _ready_fsm___pip_5160_1_124 = (_q__idx_fsm___pip_5160_1_124 == 1) || (_q__idx_fsm___pip_5160_1_124 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_124 = 0,_q__full_fsm___pip_5160_1_124 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_124 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_124 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_125,_q__idx_fsm___pip_5160_1_125;
wire _ready_fsm___pip_5160_1_125 = (_q__idx_fsm___pip_5160_1_125 == 1) || (_q__idx_fsm___pip_5160_1_125 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_125 = 0,_q__full_fsm___pip_5160_1_125 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_125 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_125 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_126,_q__idx_fsm___pip_5160_1_126;
wire _ready_fsm___pip_5160_1_126 = (_q__idx_fsm___pip_5160_1_126 == 1) || (_q__idx_fsm___pip_5160_1_126 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_126 = 0,_q__full_fsm___pip_5160_1_126 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_126 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_126 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_127,_q__idx_fsm___pip_5160_1_127;
wire _ready_fsm___pip_5160_1_127 = (_q__idx_fsm___pip_5160_1_127 == 1) || (_q__idx_fsm___pip_5160_1_127 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_127 = 0,_q__full_fsm___pip_5160_1_127 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_127 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_127 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_128,_q__idx_fsm___pip_5160_1_128;
wire _ready_fsm___pip_5160_1_128 = (_q__idx_fsm___pip_5160_1_128 == 1) || (_q__idx_fsm___pip_5160_1_128 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_128 = 0,_q__full_fsm___pip_5160_1_128 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_128 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_128 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_129,_q__idx_fsm___pip_5160_1_129;
wire _ready_fsm___pip_5160_1_129 = (_q__idx_fsm___pip_5160_1_129 == 1) || (_q__idx_fsm___pip_5160_1_129 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_129 = 0,_q__full_fsm___pip_5160_1_129 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_129 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_129 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_130,_q__idx_fsm___pip_5160_1_130;
wire _ready_fsm___pip_5160_1_130 = (_q__idx_fsm___pip_5160_1_130 == 1) || (_q__idx_fsm___pip_5160_1_130 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_130 = 0,_q__full_fsm___pip_5160_1_130 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_130 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_130 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_131,_q__idx_fsm___pip_5160_1_131;
wire _ready_fsm___pip_5160_1_131 = (_q__idx_fsm___pip_5160_1_131 == 1) || (_q__idx_fsm___pip_5160_1_131 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_131 = 0,_q__full_fsm___pip_5160_1_131 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_131 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_131 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_132,_q__idx_fsm___pip_5160_1_132;
wire _ready_fsm___pip_5160_1_132 = (_q__idx_fsm___pip_5160_1_132 == 1) || (_q__idx_fsm___pip_5160_1_132 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_132 = 0,_q__full_fsm___pip_5160_1_132 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_132 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_132 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_133,_q__idx_fsm___pip_5160_1_133;
wire _ready_fsm___pip_5160_1_133 = (_q__idx_fsm___pip_5160_1_133 == 1) || (_q__idx_fsm___pip_5160_1_133 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_133 = 0,_q__full_fsm___pip_5160_1_133 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_133 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_133 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_134,_q__idx_fsm___pip_5160_1_134;
wire _ready_fsm___pip_5160_1_134 = (_q__idx_fsm___pip_5160_1_134 == 1) || (_q__idx_fsm___pip_5160_1_134 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_134 = 0,_q__full_fsm___pip_5160_1_134 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_134 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_134 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_135,_q__idx_fsm___pip_5160_1_135;
wire _ready_fsm___pip_5160_1_135 = (_q__idx_fsm___pip_5160_1_135 == 1) || (_q__idx_fsm___pip_5160_1_135 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_135 = 0,_q__full_fsm___pip_5160_1_135 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_135 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_135 = 0;
reg  [0:0] _d__idx_fsm___pip_5160_1_136,_q__idx_fsm___pip_5160_1_136;
wire _ready_fsm___pip_5160_1_136 = (_q__idx_fsm___pip_5160_1_136 == 1) || (_q__idx_fsm___pip_5160_1_136 == 0);
reg  [0:0] _d__full_fsm___pip_5160_1_136 = 0,_q__full_fsm___pip_5160_1_136 = 0;
reg  [0:0] _t__stall_fsm___pip_5160_1_136 = 0;
reg  [0:0] _t__1stdisable_fsm___pip_5160_1_136 = 0;
assign out_pix_r = _d_pix_r;
assign out_pix_g = _d_pix_g;
assign out_pix_b = _d_pix_b;
assign out_done = (_q__idx_fsm0 == 0) && _autorun
 &&   _q__idx_fsm___pip_5160_1_0 == 0 && ~ _q__full_fsm___pip_5160_1_0
 &&   _q__idx_fsm___pip_5160_1_1 == 0 && ~ _q__full_fsm___pip_5160_1_1
 &&   _q__idx_fsm___pip_5160_1_2 == 0 && ~ _q__full_fsm___pip_5160_1_2
 &&   _q__idx_fsm___pip_5160_1_3 == 0 && ~ _q__full_fsm___pip_5160_1_3
 &&   _q__idx_fsm___pip_5160_1_4 == 0 && ~ _q__full_fsm___pip_5160_1_4
 &&   _q__idx_fsm___pip_5160_1_5 == 0 && ~ _q__full_fsm___pip_5160_1_5
 &&   _q__idx_fsm___pip_5160_1_6 == 0 && ~ _q__full_fsm___pip_5160_1_6
 &&   _q__idx_fsm___pip_5160_1_7 == 0 && ~ _q__full_fsm___pip_5160_1_7
 &&   _q__idx_fsm___pip_5160_1_8 == 0 && ~ _q__full_fsm___pip_5160_1_8
 &&   _q__idx_fsm___pip_5160_1_9 == 0 && ~ _q__full_fsm___pip_5160_1_9
 &&   _q__idx_fsm___pip_5160_1_10 == 0 && ~ _q__full_fsm___pip_5160_1_10
 &&   _q__idx_fsm___pip_5160_1_11 == 0 && ~ _q__full_fsm___pip_5160_1_11
 &&   _q__idx_fsm___pip_5160_1_12 == 0 && ~ _q__full_fsm___pip_5160_1_12
 &&   _q__idx_fsm___pip_5160_1_13 == 0 && ~ _q__full_fsm___pip_5160_1_13
 &&   _q__idx_fsm___pip_5160_1_14 == 0 && ~ _q__full_fsm___pip_5160_1_14
 &&   _q__idx_fsm___pip_5160_1_15 == 0 && ~ _q__full_fsm___pip_5160_1_15
 &&   _q__idx_fsm___pip_5160_1_16 == 0 && ~ _q__full_fsm___pip_5160_1_16
 &&   _q__idx_fsm___pip_5160_1_17 == 0 && ~ _q__full_fsm___pip_5160_1_17
 &&   _q__idx_fsm___pip_5160_1_18 == 0 && ~ _q__full_fsm___pip_5160_1_18
 &&   _q__idx_fsm___pip_5160_1_19 == 0 && ~ _q__full_fsm___pip_5160_1_19
 &&   _q__idx_fsm___pip_5160_1_20 == 0 && ~ _q__full_fsm___pip_5160_1_20
 &&   _q__idx_fsm___pip_5160_1_21 == 0 && ~ _q__full_fsm___pip_5160_1_21
 &&   _q__idx_fsm___pip_5160_1_22 == 0 && ~ _q__full_fsm___pip_5160_1_22
 &&   _q__idx_fsm___pip_5160_1_23 == 0 && ~ _q__full_fsm___pip_5160_1_23
 &&   _q__idx_fsm___pip_5160_1_24 == 0 && ~ _q__full_fsm___pip_5160_1_24
 &&   _q__idx_fsm___pip_5160_1_25 == 0 && ~ _q__full_fsm___pip_5160_1_25
 &&   _q__idx_fsm___pip_5160_1_26 == 0 && ~ _q__full_fsm___pip_5160_1_26
 &&   _q__idx_fsm___pip_5160_1_27 == 0 && ~ _q__full_fsm___pip_5160_1_27
 &&   _q__idx_fsm___pip_5160_1_28 == 0 && ~ _q__full_fsm___pip_5160_1_28
 &&   _q__idx_fsm___pip_5160_1_29 == 0 && ~ _q__full_fsm___pip_5160_1_29
 &&   _q__idx_fsm___pip_5160_1_30 == 0 && ~ _q__full_fsm___pip_5160_1_30
 &&   _q__idx_fsm___pip_5160_1_31 == 0 && ~ _q__full_fsm___pip_5160_1_31
 &&   _q__idx_fsm___pip_5160_1_32 == 0 && ~ _q__full_fsm___pip_5160_1_32
 &&   _q__idx_fsm___pip_5160_1_33 == 0 && ~ _q__full_fsm___pip_5160_1_33
 &&   _q__idx_fsm___pip_5160_1_34 == 0 && ~ _q__full_fsm___pip_5160_1_34
 &&   _q__idx_fsm___pip_5160_1_35 == 0 && ~ _q__full_fsm___pip_5160_1_35
 &&   _q__idx_fsm___pip_5160_1_36 == 0 && ~ _q__full_fsm___pip_5160_1_36
 &&   _q__idx_fsm___pip_5160_1_37 == 0 && ~ _q__full_fsm___pip_5160_1_37
 &&   _q__idx_fsm___pip_5160_1_38 == 0 && ~ _q__full_fsm___pip_5160_1_38
 &&   _q__idx_fsm___pip_5160_1_39 == 0 && ~ _q__full_fsm___pip_5160_1_39
 &&   _q__idx_fsm___pip_5160_1_40 == 0 && ~ _q__full_fsm___pip_5160_1_40
 &&   _q__idx_fsm___pip_5160_1_41 == 0 && ~ _q__full_fsm___pip_5160_1_41
 &&   _q__idx_fsm___pip_5160_1_42 == 0 && ~ _q__full_fsm___pip_5160_1_42
 &&   _q__idx_fsm___pip_5160_1_43 == 0 && ~ _q__full_fsm___pip_5160_1_43
 &&   _q__idx_fsm___pip_5160_1_44 == 0 && ~ _q__full_fsm___pip_5160_1_44
 &&   _q__idx_fsm___pip_5160_1_45 == 0 && ~ _q__full_fsm___pip_5160_1_45
 &&   _q__idx_fsm___pip_5160_1_46 == 0 && ~ _q__full_fsm___pip_5160_1_46
 &&   _q__idx_fsm___pip_5160_1_47 == 0 && ~ _q__full_fsm___pip_5160_1_47
 &&   _q__idx_fsm___pip_5160_1_48 == 0 && ~ _q__full_fsm___pip_5160_1_48
 &&   _q__idx_fsm___pip_5160_1_49 == 0 && ~ _q__full_fsm___pip_5160_1_49
 &&   _q__idx_fsm___pip_5160_1_50 == 0 && ~ _q__full_fsm___pip_5160_1_50
 &&   _q__idx_fsm___pip_5160_1_51 == 0 && ~ _q__full_fsm___pip_5160_1_51
 &&   _q__idx_fsm___pip_5160_1_52 == 0 && ~ _q__full_fsm___pip_5160_1_52
 &&   _q__idx_fsm___pip_5160_1_53 == 0 && ~ _q__full_fsm___pip_5160_1_53
 &&   _q__idx_fsm___pip_5160_1_54 == 0 && ~ _q__full_fsm___pip_5160_1_54
 &&   _q__idx_fsm___pip_5160_1_55 == 0 && ~ _q__full_fsm___pip_5160_1_55
 &&   _q__idx_fsm___pip_5160_1_56 == 0 && ~ _q__full_fsm___pip_5160_1_56
 &&   _q__idx_fsm___pip_5160_1_57 == 0 && ~ _q__full_fsm___pip_5160_1_57
 &&   _q__idx_fsm___pip_5160_1_58 == 0 && ~ _q__full_fsm___pip_5160_1_58
 &&   _q__idx_fsm___pip_5160_1_59 == 0 && ~ _q__full_fsm___pip_5160_1_59
 &&   _q__idx_fsm___pip_5160_1_60 == 0 && ~ _q__full_fsm___pip_5160_1_60
 &&   _q__idx_fsm___pip_5160_1_61 == 0 && ~ _q__full_fsm___pip_5160_1_61
 &&   _q__idx_fsm___pip_5160_1_62 == 0 && ~ _q__full_fsm___pip_5160_1_62
 &&   _q__idx_fsm___pip_5160_1_63 == 0 && ~ _q__full_fsm___pip_5160_1_63
 &&   _q__idx_fsm___pip_5160_1_64 == 0 && ~ _q__full_fsm___pip_5160_1_64
 &&   _q__idx_fsm___pip_5160_1_65 == 0 && ~ _q__full_fsm___pip_5160_1_65
 &&   _q__idx_fsm___pip_5160_1_66 == 0 && ~ _q__full_fsm___pip_5160_1_66
 &&   _q__idx_fsm___pip_5160_1_67 == 0 && ~ _q__full_fsm___pip_5160_1_67
 &&   _q__idx_fsm___pip_5160_1_68 == 0 && ~ _q__full_fsm___pip_5160_1_68
 &&   _q__idx_fsm___pip_5160_1_69 == 0 && ~ _q__full_fsm___pip_5160_1_69
 &&   _q__idx_fsm___pip_5160_1_70 == 0 && ~ _q__full_fsm___pip_5160_1_70
 &&   _q__idx_fsm___pip_5160_1_71 == 0 && ~ _q__full_fsm___pip_5160_1_71
 &&   _q__idx_fsm___pip_5160_1_72 == 0 && ~ _q__full_fsm___pip_5160_1_72
 &&   _q__idx_fsm___pip_5160_1_73 == 0 && ~ _q__full_fsm___pip_5160_1_73
 &&   _q__idx_fsm___pip_5160_1_74 == 0 && ~ _q__full_fsm___pip_5160_1_74
 &&   _q__idx_fsm___pip_5160_1_75 == 0 && ~ _q__full_fsm___pip_5160_1_75
 &&   _q__idx_fsm___pip_5160_1_76 == 0 && ~ _q__full_fsm___pip_5160_1_76
 &&   _q__idx_fsm___pip_5160_1_77 == 0 && ~ _q__full_fsm___pip_5160_1_77
 &&   _q__idx_fsm___pip_5160_1_78 == 0 && ~ _q__full_fsm___pip_5160_1_78
 &&   _q__idx_fsm___pip_5160_1_79 == 0 && ~ _q__full_fsm___pip_5160_1_79
 &&   _q__idx_fsm___pip_5160_1_80 == 0 && ~ _q__full_fsm___pip_5160_1_80
 &&   _q__idx_fsm___pip_5160_1_81 == 0 && ~ _q__full_fsm___pip_5160_1_81
 &&   _q__idx_fsm___pip_5160_1_82 == 0 && ~ _q__full_fsm___pip_5160_1_82
 &&   _q__idx_fsm___pip_5160_1_83 == 0 && ~ _q__full_fsm___pip_5160_1_83
 &&   _q__idx_fsm___pip_5160_1_84 == 0 && ~ _q__full_fsm___pip_5160_1_84
 &&   _q__idx_fsm___pip_5160_1_85 == 0 && ~ _q__full_fsm___pip_5160_1_85
 &&   _q__idx_fsm___pip_5160_1_86 == 0 && ~ _q__full_fsm___pip_5160_1_86
 &&   _q__idx_fsm___pip_5160_1_87 == 0 && ~ _q__full_fsm___pip_5160_1_87
 &&   _q__idx_fsm___pip_5160_1_88 == 0 && ~ _q__full_fsm___pip_5160_1_88
 &&   _q__idx_fsm___pip_5160_1_89 == 0 && ~ _q__full_fsm___pip_5160_1_89
 &&   _q__idx_fsm___pip_5160_1_90 == 0 && ~ _q__full_fsm___pip_5160_1_90
 &&   _q__idx_fsm___pip_5160_1_91 == 0 && ~ _q__full_fsm___pip_5160_1_91
 &&   _q__idx_fsm___pip_5160_1_92 == 0 && ~ _q__full_fsm___pip_5160_1_92
 &&   _q__idx_fsm___pip_5160_1_93 == 0 && ~ _q__full_fsm___pip_5160_1_93
 &&   _q__idx_fsm___pip_5160_1_94 == 0 && ~ _q__full_fsm___pip_5160_1_94
 &&   _q__idx_fsm___pip_5160_1_95 == 0 && ~ _q__full_fsm___pip_5160_1_95
 &&   _q__idx_fsm___pip_5160_1_96 == 0 && ~ _q__full_fsm___pip_5160_1_96
 &&   _q__idx_fsm___pip_5160_1_97 == 0 && ~ _q__full_fsm___pip_5160_1_97
 &&   _q__idx_fsm___pip_5160_1_98 == 0 && ~ _q__full_fsm___pip_5160_1_98
 &&   _q__idx_fsm___pip_5160_1_99 == 0 && ~ _q__full_fsm___pip_5160_1_99
 &&   _q__idx_fsm___pip_5160_1_100 == 0 && ~ _q__full_fsm___pip_5160_1_100
 &&   _q__idx_fsm___pip_5160_1_101 == 0 && ~ _q__full_fsm___pip_5160_1_101
 &&   _q__idx_fsm___pip_5160_1_102 == 0 && ~ _q__full_fsm___pip_5160_1_102
 &&   _q__idx_fsm___pip_5160_1_103 == 0 && ~ _q__full_fsm___pip_5160_1_103
 &&   _q__idx_fsm___pip_5160_1_104 == 0 && ~ _q__full_fsm___pip_5160_1_104
 &&   _q__idx_fsm___pip_5160_1_105 == 0 && ~ _q__full_fsm___pip_5160_1_105
 &&   _q__idx_fsm___pip_5160_1_106 == 0 && ~ _q__full_fsm___pip_5160_1_106
 &&   _q__idx_fsm___pip_5160_1_107 == 0 && ~ _q__full_fsm___pip_5160_1_107
 &&   _q__idx_fsm___pip_5160_1_108 == 0 && ~ _q__full_fsm___pip_5160_1_108
 &&   _q__idx_fsm___pip_5160_1_109 == 0 && ~ _q__full_fsm___pip_5160_1_109
 &&   _q__idx_fsm___pip_5160_1_110 == 0 && ~ _q__full_fsm___pip_5160_1_110
 &&   _q__idx_fsm___pip_5160_1_111 == 0 && ~ _q__full_fsm___pip_5160_1_111
 &&   _q__idx_fsm___pip_5160_1_112 == 0 && ~ _q__full_fsm___pip_5160_1_112
 &&   _q__idx_fsm___pip_5160_1_113 == 0 && ~ _q__full_fsm___pip_5160_1_113
 &&   _q__idx_fsm___pip_5160_1_114 == 0 && ~ _q__full_fsm___pip_5160_1_114
 &&   _q__idx_fsm___pip_5160_1_115 == 0 && ~ _q__full_fsm___pip_5160_1_115
 &&   _q__idx_fsm___pip_5160_1_116 == 0 && ~ _q__full_fsm___pip_5160_1_116
 &&   _q__idx_fsm___pip_5160_1_117 == 0 && ~ _q__full_fsm___pip_5160_1_117
 &&   _q__idx_fsm___pip_5160_1_118 == 0 && ~ _q__full_fsm___pip_5160_1_118
 &&   _q__idx_fsm___pip_5160_1_119 == 0 && ~ _q__full_fsm___pip_5160_1_119
 &&   _q__idx_fsm___pip_5160_1_120 == 0 && ~ _q__full_fsm___pip_5160_1_120
 &&   _q__idx_fsm___pip_5160_1_121 == 0 && ~ _q__full_fsm___pip_5160_1_121
 &&   _q__idx_fsm___pip_5160_1_122 == 0 && ~ _q__full_fsm___pip_5160_1_122
 &&   _q__idx_fsm___pip_5160_1_123 == 0 && ~ _q__full_fsm___pip_5160_1_123
 &&   _q__idx_fsm___pip_5160_1_124 == 0 && ~ _q__full_fsm___pip_5160_1_124
 &&   _q__idx_fsm___pip_5160_1_125 == 0 && ~ _q__full_fsm___pip_5160_1_125
 &&   _q__idx_fsm___pip_5160_1_126 == 0 && ~ _q__full_fsm___pip_5160_1_126
 &&   _q__idx_fsm___pip_5160_1_127 == 0 && ~ _q__full_fsm___pip_5160_1_127
 &&   _q__idx_fsm___pip_5160_1_128 == 0 && ~ _q__full_fsm___pip_5160_1_128
 &&   _q__idx_fsm___pip_5160_1_129 == 0 && ~ _q__full_fsm___pip_5160_1_129
 &&   _q__idx_fsm___pip_5160_1_130 == 0 && ~ _q__full_fsm___pip_5160_1_130
 &&   _q__idx_fsm___pip_5160_1_131 == 0 && ~ _q__full_fsm___pip_5160_1_131
 &&   _q__idx_fsm___pip_5160_1_132 == 0 && ~ _q__full_fsm___pip_5160_1_132
 &&   _q__idx_fsm___pip_5160_1_133 == 0 && ~ _q__full_fsm___pip_5160_1_133
 &&   _q__idx_fsm___pip_5160_1_134 == 0 && ~ _q__full_fsm___pip_5160_1_134
 &&   _q__idx_fsm___pip_5160_1_135 == 0 && ~ _q__full_fsm___pip_5160_1_135
 &&   _q__idx_fsm___pip_5160_1_136 == 0
;

M_frame_display__mem_cos __mem__cos(
.clock0(clock),
.clock1(clock),
.in_wenable0(_t_cos_wenable0),
.in_wdata0(_t_cos_wdata0),
.in_addr0(_d_cos_addr0),
.in_wenable1(_t_cos_wenable1),
.in_wdata1(_t_cos_wdata1),
.in_addr1(_d_cos_addr1),
.out_rdata0(_w_mem_cos_rdata0),
.out_rdata1(_w_mem_cos_rdata1)
);
M_frame_display__mem_sin __mem__sin(
.clock0(clock),
.clock1(clock),
.in_wenable0(_t_sin_wenable0),
.in_wdata0(_t_sin_wdata0),
.in_addr0(_d_sin_addr0),
.in_wenable1(_t_sin_wenable1),
.in_wdata1(_t_sin_wdata1),
.in_addr1(_d_sin_addr1),
.out_rdata0(_w_mem_sin_rdata0),
.out_rdata1(_w_mem_sin_rdata1)
);
M_frame_display__mem_invA __mem__invA(
.clock0(clock),
.clock1(clock),
.in_wenable0(_t_invA_wenable0),
.in_wdata0(_t_invA_wdata0),
.in_addr0(_d_invA_addr0),
.in_wenable1(_t_invA_wenable1),
.in_wdata1(_t_invA_wdata1),
.in_addr1(_d_invA_addr1),
.out_rdata0(_w_mem_invA_rdata0),
.out_rdata1(_w_mem_invA_rdata1)
);
M_frame_display__mem_invB __mem__invB(
.clock(clock),
.in_wenable(_t_invB_wenable),
.in_wdata(_t_invB_wdata),
.in_addr(_d_invB_addr),
.out_rdata(_w_mem_invB_rdata)
);

assign _w_tile = {1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1};

`ifdef FORMAL
initial begin
assume(reset);
end
assume property($initstate || (out_done));
`endif
always @* begin
_d_frame = _q_frame;
_d_cos_addr0 = _q_cos_addr0;
_d_cos_addr1 = _q_cos_addr1;
_d_sin_addr0 = _q_sin_addr0;
_d_sin_addr1 = _q_sin_addr1;
_d_invA_addr0 = _q_invA_addr0;
_d_invA_addr1 = _q_invA_addr1;
_d_invB_addr = _q_invB_addr;
_d___pip_5160_1_3___block_25_r_x_delta = _q___pip_5160_1_3___block_25_r_x_delta;
_d___pip_5160_1_4___block_25_r_x_delta = _q___pip_5160_1_4___block_25_r_x_delta;
_d___pip_5160_1_3___block_25_r_z_delta = _q___pip_5160_1_3___block_25_r_z_delta;
_d___pip_5160_1_4___block_25_r_z_delta = _q___pip_5160_1_4___block_25_r_z_delta;
_d___pip_5160_1_135___block_2731_clr_b = _q___pip_5160_1_135___block_2731_clr_b;
_d___pip_5160_1_136___block_2731_clr_b = _q___pip_5160_1_136___block_2731_clr_b;
_d___pip_5160_1_135___block_2731_clr_g = _q___pip_5160_1_135___block_2731_clr_g;
_d___pip_5160_1_136___block_2731_clr_g = _q___pip_5160_1_136___block_2731_clr_g;
_d___pip_5160_1_135___block_2731_clr_r = _q___pip_5160_1_135___block_2731_clr_r;
_d___pip_5160_1_136___block_2731_clr_r = _q___pip_5160_1_136___block_2731_clr_r;
_d___pip_5160_1_6___block_34_tm_x = _q___pip_5160_1_6___block_34_tm_x;
_d___pip_5160_1_7___block_34_tm_x = _q___pip_5160_1_7___block_34_tm_x;
_d___pip_5160_1_8___block_34_tm_x = _q___pip_5160_1_8___block_34_tm_x;
_d___pip_5160_1_9___block_34_tm_x = _q___pip_5160_1_9___block_34_tm_x;
_d___pip_5160_1_10___block_34_tm_x = _q___pip_5160_1_10___block_34_tm_x;
_d___pip_5160_1_11___block_34_tm_x = _q___pip_5160_1_11___block_34_tm_x;
_d___pip_5160_1_12___block_34_tm_x = _q___pip_5160_1_12___block_34_tm_x;
_d___pip_5160_1_13___block_34_tm_x = _q___pip_5160_1_13___block_34_tm_x;
_d___pip_5160_1_14___block_34_tm_x = _q___pip_5160_1_14___block_34_tm_x;
_d___pip_5160_1_15___block_34_tm_x = _q___pip_5160_1_15___block_34_tm_x;
_d___pip_5160_1_16___block_34_tm_x = _q___pip_5160_1_16___block_34_tm_x;
_d___pip_5160_1_17___block_34_tm_x = _q___pip_5160_1_17___block_34_tm_x;
_d___pip_5160_1_18___block_34_tm_x = _q___pip_5160_1_18___block_34_tm_x;
_d___pip_5160_1_19___block_34_tm_x = _q___pip_5160_1_19___block_34_tm_x;
_d___pip_5160_1_20___block_34_tm_x = _q___pip_5160_1_20___block_34_tm_x;
_d___pip_5160_1_21___block_34_tm_x = _q___pip_5160_1_21___block_34_tm_x;
_d___pip_5160_1_22___block_34_tm_x = _q___pip_5160_1_22___block_34_tm_x;
_d___pip_5160_1_23___block_34_tm_x = _q___pip_5160_1_23___block_34_tm_x;
_d___pip_5160_1_24___block_34_tm_x = _q___pip_5160_1_24___block_34_tm_x;
_d___pip_5160_1_25___block_34_tm_x = _q___pip_5160_1_25___block_34_tm_x;
_d___pip_5160_1_26___block_34_tm_x = _q___pip_5160_1_26___block_34_tm_x;
_d___pip_5160_1_27___block_34_tm_x = _q___pip_5160_1_27___block_34_tm_x;
_d___pip_5160_1_28___block_34_tm_x = _q___pip_5160_1_28___block_34_tm_x;
_d___pip_5160_1_29___block_34_tm_x = _q___pip_5160_1_29___block_34_tm_x;
_d___pip_5160_1_30___block_34_tm_x = _q___pip_5160_1_30___block_34_tm_x;
_d___pip_5160_1_31___block_34_tm_x = _q___pip_5160_1_31___block_34_tm_x;
_d___pip_5160_1_32___block_34_tm_x = _q___pip_5160_1_32___block_34_tm_x;
_d___pip_5160_1_33___block_34_tm_x = _q___pip_5160_1_33___block_34_tm_x;
_d___pip_5160_1_34___block_34_tm_x = _q___pip_5160_1_34___block_34_tm_x;
_d___pip_5160_1_35___block_34_tm_x = _q___pip_5160_1_35___block_34_tm_x;
_d___pip_5160_1_36___block_34_tm_x = _q___pip_5160_1_36___block_34_tm_x;
_d___pip_5160_1_37___block_34_tm_x = _q___pip_5160_1_37___block_34_tm_x;
_d___pip_5160_1_38___block_34_tm_x = _q___pip_5160_1_38___block_34_tm_x;
_d___pip_5160_1_39___block_34_tm_x = _q___pip_5160_1_39___block_34_tm_x;
_d___pip_5160_1_40___block_34_tm_x = _q___pip_5160_1_40___block_34_tm_x;
_d___pip_5160_1_41___block_34_tm_x = _q___pip_5160_1_41___block_34_tm_x;
_d___pip_5160_1_42___block_34_tm_x = _q___pip_5160_1_42___block_34_tm_x;
_d___pip_5160_1_43___block_34_tm_x = _q___pip_5160_1_43___block_34_tm_x;
_d___pip_5160_1_44___block_34_tm_x = _q___pip_5160_1_44___block_34_tm_x;
_d___pip_5160_1_45___block_34_tm_x = _q___pip_5160_1_45___block_34_tm_x;
_d___pip_5160_1_46___block_34_tm_x = _q___pip_5160_1_46___block_34_tm_x;
_d___pip_5160_1_47___block_34_tm_x = _q___pip_5160_1_47___block_34_tm_x;
_d___pip_5160_1_48___block_34_tm_x = _q___pip_5160_1_48___block_34_tm_x;
_d___pip_5160_1_49___block_34_tm_x = _q___pip_5160_1_49___block_34_tm_x;
_d___pip_5160_1_50___block_34_tm_x = _q___pip_5160_1_50___block_34_tm_x;
_d___pip_5160_1_51___block_34_tm_x = _q___pip_5160_1_51___block_34_tm_x;
_d___pip_5160_1_52___block_34_tm_x = _q___pip_5160_1_52___block_34_tm_x;
_d___pip_5160_1_53___block_34_tm_x = _q___pip_5160_1_53___block_34_tm_x;
_d___pip_5160_1_54___block_34_tm_x = _q___pip_5160_1_54___block_34_tm_x;
_d___pip_5160_1_55___block_34_tm_x = _q___pip_5160_1_55___block_34_tm_x;
_d___pip_5160_1_56___block_34_tm_x = _q___pip_5160_1_56___block_34_tm_x;
_d___pip_5160_1_57___block_34_tm_x = _q___pip_5160_1_57___block_34_tm_x;
_d___pip_5160_1_58___block_34_tm_x = _q___pip_5160_1_58___block_34_tm_x;
_d___pip_5160_1_59___block_34_tm_x = _q___pip_5160_1_59___block_34_tm_x;
_d___pip_5160_1_60___block_34_tm_x = _q___pip_5160_1_60___block_34_tm_x;
_d___pip_5160_1_61___block_34_tm_x = _q___pip_5160_1_61___block_34_tm_x;
_d___pip_5160_1_62___block_34_tm_x = _q___pip_5160_1_62___block_34_tm_x;
_d___pip_5160_1_63___block_34_tm_x = _q___pip_5160_1_63___block_34_tm_x;
_d___pip_5160_1_64___block_34_tm_x = _q___pip_5160_1_64___block_34_tm_x;
_d___pip_5160_1_65___block_34_tm_x = _q___pip_5160_1_65___block_34_tm_x;
_d___pip_5160_1_66___block_34_tm_x = _q___pip_5160_1_66___block_34_tm_x;
_d___pip_5160_1_67___block_34_tm_x = _q___pip_5160_1_67___block_34_tm_x;
_d___pip_5160_1_68___block_34_tm_x = _q___pip_5160_1_68___block_34_tm_x;
_d___pip_5160_1_69___block_34_tm_x = _q___pip_5160_1_69___block_34_tm_x;
_d___pip_5160_1_70___block_34_tm_x = _q___pip_5160_1_70___block_34_tm_x;
_d___pip_5160_1_71___block_34_tm_x = _q___pip_5160_1_71___block_34_tm_x;
_d___pip_5160_1_72___block_34_tm_x = _q___pip_5160_1_72___block_34_tm_x;
_d___pip_5160_1_73___block_34_tm_x = _q___pip_5160_1_73___block_34_tm_x;
_d___pip_5160_1_74___block_34_tm_x = _q___pip_5160_1_74___block_34_tm_x;
_d___pip_5160_1_75___block_34_tm_x = _q___pip_5160_1_75___block_34_tm_x;
_d___pip_5160_1_76___block_34_tm_x = _q___pip_5160_1_76___block_34_tm_x;
_d___pip_5160_1_77___block_34_tm_x = _q___pip_5160_1_77___block_34_tm_x;
_d___pip_5160_1_78___block_34_tm_x = _q___pip_5160_1_78___block_34_tm_x;
_d___pip_5160_1_79___block_34_tm_x = _q___pip_5160_1_79___block_34_tm_x;
_d___pip_5160_1_80___block_34_tm_x = _q___pip_5160_1_80___block_34_tm_x;
_d___pip_5160_1_81___block_34_tm_x = _q___pip_5160_1_81___block_34_tm_x;
_d___pip_5160_1_82___block_34_tm_x = _q___pip_5160_1_82___block_34_tm_x;
_d___pip_5160_1_83___block_34_tm_x = _q___pip_5160_1_83___block_34_tm_x;
_d___pip_5160_1_84___block_34_tm_x = _q___pip_5160_1_84___block_34_tm_x;
_d___pip_5160_1_85___block_34_tm_x = _q___pip_5160_1_85___block_34_tm_x;
_d___pip_5160_1_86___block_34_tm_x = _q___pip_5160_1_86___block_34_tm_x;
_d___pip_5160_1_87___block_34_tm_x = _q___pip_5160_1_87___block_34_tm_x;
_d___pip_5160_1_88___block_34_tm_x = _q___pip_5160_1_88___block_34_tm_x;
_d___pip_5160_1_89___block_34_tm_x = _q___pip_5160_1_89___block_34_tm_x;
_d___pip_5160_1_90___block_34_tm_x = _q___pip_5160_1_90___block_34_tm_x;
_d___pip_5160_1_91___block_34_tm_x = _q___pip_5160_1_91___block_34_tm_x;
_d___pip_5160_1_92___block_34_tm_x = _q___pip_5160_1_92___block_34_tm_x;
_d___pip_5160_1_93___block_34_tm_x = _q___pip_5160_1_93___block_34_tm_x;
_d___pip_5160_1_94___block_34_tm_x = _q___pip_5160_1_94___block_34_tm_x;
_d___pip_5160_1_95___block_34_tm_x = _q___pip_5160_1_95___block_34_tm_x;
_d___pip_5160_1_96___block_34_tm_x = _q___pip_5160_1_96___block_34_tm_x;
_d___pip_5160_1_97___block_34_tm_x = _q___pip_5160_1_97___block_34_tm_x;
_d___pip_5160_1_98___block_34_tm_x = _q___pip_5160_1_98___block_34_tm_x;
_d___pip_5160_1_99___block_34_tm_x = _q___pip_5160_1_99___block_34_tm_x;
_d___pip_5160_1_100___block_34_tm_x = _q___pip_5160_1_100___block_34_tm_x;
_d___pip_5160_1_101___block_34_tm_x = _q___pip_5160_1_101___block_34_tm_x;
_d___pip_5160_1_102___block_34_tm_x = _q___pip_5160_1_102___block_34_tm_x;
_d___pip_5160_1_103___block_34_tm_x = _q___pip_5160_1_103___block_34_tm_x;
_d___pip_5160_1_104___block_34_tm_x = _q___pip_5160_1_104___block_34_tm_x;
_d___pip_5160_1_105___block_34_tm_x = _q___pip_5160_1_105___block_34_tm_x;
_d___pip_5160_1_106___block_34_tm_x = _q___pip_5160_1_106___block_34_tm_x;
_d___pip_5160_1_107___block_34_tm_x = _q___pip_5160_1_107___block_34_tm_x;
_d___pip_5160_1_108___block_34_tm_x = _q___pip_5160_1_108___block_34_tm_x;
_d___pip_5160_1_109___block_34_tm_x = _q___pip_5160_1_109___block_34_tm_x;
_d___pip_5160_1_110___block_34_tm_x = _q___pip_5160_1_110___block_34_tm_x;
_d___pip_5160_1_111___block_34_tm_x = _q___pip_5160_1_111___block_34_tm_x;
_d___pip_5160_1_112___block_34_tm_x = _q___pip_5160_1_112___block_34_tm_x;
_d___pip_5160_1_113___block_34_tm_x = _q___pip_5160_1_113___block_34_tm_x;
_d___pip_5160_1_114___block_34_tm_x = _q___pip_5160_1_114___block_34_tm_x;
_d___pip_5160_1_115___block_34_tm_x = _q___pip_5160_1_115___block_34_tm_x;
_d___pip_5160_1_116___block_34_tm_x = _q___pip_5160_1_116___block_34_tm_x;
_d___pip_5160_1_117___block_34_tm_x = _q___pip_5160_1_117___block_34_tm_x;
_d___pip_5160_1_118___block_34_tm_x = _q___pip_5160_1_118___block_34_tm_x;
_d___pip_5160_1_119___block_34_tm_x = _q___pip_5160_1_119___block_34_tm_x;
_d___pip_5160_1_120___block_34_tm_x = _q___pip_5160_1_120___block_34_tm_x;
_d___pip_5160_1_121___block_34_tm_x = _q___pip_5160_1_121___block_34_tm_x;
_d___pip_5160_1_122___block_34_tm_x = _q___pip_5160_1_122___block_34_tm_x;
_d___pip_5160_1_123___block_34_tm_x = _q___pip_5160_1_123___block_34_tm_x;
_d___pip_5160_1_124___block_34_tm_x = _q___pip_5160_1_124___block_34_tm_x;
_d___pip_5160_1_125___block_34_tm_x = _q___pip_5160_1_125___block_34_tm_x;
_d___pip_5160_1_126___block_34_tm_x = _q___pip_5160_1_126___block_34_tm_x;
_d___pip_5160_1_127___block_34_tm_x = _q___pip_5160_1_127___block_34_tm_x;
_d___pip_5160_1_128___block_34_tm_x = _q___pip_5160_1_128___block_34_tm_x;
_d___pip_5160_1_129___block_34_tm_x = _q___pip_5160_1_129___block_34_tm_x;
_d___pip_5160_1_130___block_34_tm_x = _q___pip_5160_1_130___block_34_tm_x;
_d___pip_5160_1_131___block_34_tm_x = _q___pip_5160_1_131___block_34_tm_x;
_d___pip_5160_1_132___block_34_tm_x = _q___pip_5160_1_132___block_34_tm_x;
_d___pip_5160_1_133___block_34_tm_x = _q___pip_5160_1_133___block_34_tm_x;
_d___pip_5160_1_134___block_34_tm_x = _q___pip_5160_1_134___block_34_tm_x;
_d___pip_5160_1_6___block_34_tm_y = _q___pip_5160_1_6___block_34_tm_y;
_d___pip_5160_1_7___block_34_tm_y = _q___pip_5160_1_7___block_34_tm_y;
_d___pip_5160_1_8___block_34_tm_y = _q___pip_5160_1_8___block_34_tm_y;
_d___pip_5160_1_9___block_34_tm_y = _q___pip_5160_1_9___block_34_tm_y;
_d___pip_5160_1_10___block_34_tm_y = _q___pip_5160_1_10___block_34_tm_y;
_d___pip_5160_1_11___block_34_tm_y = _q___pip_5160_1_11___block_34_tm_y;
_d___pip_5160_1_12___block_34_tm_y = _q___pip_5160_1_12___block_34_tm_y;
_d___pip_5160_1_13___block_34_tm_y = _q___pip_5160_1_13___block_34_tm_y;
_d___pip_5160_1_14___block_34_tm_y = _q___pip_5160_1_14___block_34_tm_y;
_d___pip_5160_1_15___block_34_tm_y = _q___pip_5160_1_15___block_34_tm_y;
_d___pip_5160_1_16___block_34_tm_y = _q___pip_5160_1_16___block_34_tm_y;
_d___pip_5160_1_17___block_34_tm_y = _q___pip_5160_1_17___block_34_tm_y;
_d___pip_5160_1_18___block_34_tm_y = _q___pip_5160_1_18___block_34_tm_y;
_d___pip_5160_1_19___block_34_tm_y = _q___pip_5160_1_19___block_34_tm_y;
_d___pip_5160_1_20___block_34_tm_y = _q___pip_5160_1_20___block_34_tm_y;
_d___pip_5160_1_21___block_34_tm_y = _q___pip_5160_1_21___block_34_tm_y;
_d___pip_5160_1_22___block_34_tm_y = _q___pip_5160_1_22___block_34_tm_y;
_d___pip_5160_1_23___block_34_tm_y = _q___pip_5160_1_23___block_34_tm_y;
_d___pip_5160_1_24___block_34_tm_y = _q___pip_5160_1_24___block_34_tm_y;
_d___pip_5160_1_25___block_34_tm_y = _q___pip_5160_1_25___block_34_tm_y;
_d___pip_5160_1_26___block_34_tm_y = _q___pip_5160_1_26___block_34_tm_y;
_d___pip_5160_1_27___block_34_tm_y = _q___pip_5160_1_27___block_34_tm_y;
_d___pip_5160_1_28___block_34_tm_y = _q___pip_5160_1_28___block_34_tm_y;
_d___pip_5160_1_29___block_34_tm_y = _q___pip_5160_1_29___block_34_tm_y;
_d___pip_5160_1_30___block_34_tm_y = _q___pip_5160_1_30___block_34_tm_y;
_d___pip_5160_1_31___block_34_tm_y = _q___pip_5160_1_31___block_34_tm_y;
_d___pip_5160_1_32___block_34_tm_y = _q___pip_5160_1_32___block_34_tm_y;
_d___pip_5160_1_33___block_34_tm_y = _q___pip_5160_1_33___block_34_tm_y;
_d___pip_5160_1_34___block_34_tm_y = _q___pip_5160_1_34___block_34_tm_y;
_d___pip_5160_1_35___block_34_tm_y = _q___pip_5160_1_35___block_34_tm_y;
_d___pip_5160_1_36___block_34_tm_y = _q___pip_5160_1_36___block_34_tm_y;
_d___pip_5160_1_37___block_34_tm_y = _q___pip_5160_1_37___block_34_tm_y;
_d___pip_5160_1_38___block_34_tm_y = _q___pip_5160_1_38___block_34_tm_y;
_d___pip_5160_1_39___block_34_tm_y = _q___pip_5160_1_39___block_34_tm_y;
_d___pip_5160_1_40___block_34_tm_y = _q___pip_5160_1_40___block_34_tm_y;
_d___pip_5160_1_41___block_34_tm_y = _q___pip_5160_1_41___block_34_tm_y;
_d___pip_5160_1_42___block_34_tm_y = _q___pip_5160_1_42___block_34_tm_y;
_d___pip_5160_1_43___block_34_tm_y = _q___pip_5160_1_43___block_34_tm_y;
_d___pip_5160_1_44___block_34_tm_y = _q___pip_5160_1_44___block_34_tm_y;
_d___pip_5160_1_45___block_34_tm_y = _q___pip_5160_1_45___block_34_tm_y;
_d___pip_5160_1_46___block_34_tm_y = _q___pip_5160_1_46___block_34_tm_y;
_d___pip_5160_1_47___block_34_tm_y = _q___pip_5160_1_47___block_34_tm_y;
_d___pip_5160_1_48___block_34_tm_y = _q___pip_5160_1_48___block_34_tm_y;
_d___pip_5160_1_49___block_34_tm_y = _q___pip_5160_1_49___block_34_tm_y;
_d___pip_5160_1_50___block_34_tm_y = _q___pip_5160_1_50___block_34_tm_y;
_d___pip_5160_1_51___block_34_tm_y = _q___pip_5160_1_51___block_34_tm_y;
_d___pip_5160_1_52___block_34_tm_y = _q___pip_5160_1_52___block_34_tm_y;
_d___pip_5160_1_53___block_34_tm_y = _q___pip_5160_1_53___block_34_tm_y;
_d___pip_5160_1_54___block_34_tm_y = _q___pip_5160_1_54___block_34_tm_y;
_d___pip_5160_1_55___block_34_tm_y = _q___pip_5160_1_55___block_34_tm_y;
_d___pip_5160_1_56___block_34_tm_y = _q___pip_5160_1_56___block_34_tm_y;
_d___pip_5160_1_57___block_34_tm_y = _q___pip_5160_1_57___block_34_tm_y;
_d___pip_5160_1_58___block_34_tm_y = _q___pip_5160_1_58___block_34_tm_y;
_d___pip_5160_1_59___block_34_tm_y = _q___pip_5160_1_59___block_34_tm_y;
_d___pip_5160_1_60___block_34_tm_y = _q___pip_5160_1_60___block_34_tm_y;
_d___pip_5160_1_61___block_34_tm_y = _q___pip_5160_1_61___block_34_tm_y;
_d___pip_5160_1_62___block_34_tm_y = _q___pip_5160_1_62___block_34_tm_y;
_d___pip_5160_1_63___block_34_tm_y = _q___pip_5160_1_63___block_34_tm_y;
_d___pip_5160_1_64___block_34_tm_y = _q___pip_5160_1_64___block_34_tm_y;
_d___pip_5160_1_65___block_34_tm_y = _q___pip_5160_1_65___block_34_tm_y;
_d___pip_5160_1_66___block_34_tm_y = _q___pip_5160_1_66___block_34_tm_y;
_d___pip_5160_1_67___block_34_tm_y = _q___pip_5160_1_67___block_34_tm_y;
_d___pip_5160_1_68___block_34_tm_y = _q___pip_5160_1_68___block_34_tm_y;
_d___pip_5160_1_69___block_34_tm_y = _q___pip_5160_1_69___block_34_tm_y;
_d___pip_5160_1_70___block_34_tm_y = _q___pip_5160_1_70___block_34_tm_y;
_d___pip_5160_1_71___block_34_tm_y = _q___pip_5160_1_71___block_34_tm_y;
_d___pip_5160_1_72___block_34_tm_y = _q___pip_5160_1_72___block_34_tm_y;
_d___pip_5160_1_73___block_34_tm_y = _q___pip_5160_1_73___block_34_tm_y;
_d___pip_5160_1_74___block_34_tm_y = _q___pip_5160_1_74___block_34_tm_y;
_d___pip_5160_1_75___block_34_tm_y = _q___pip_5160_1_75___block_34_tm_y;
_d___pip_5160_1_76___block_34_tm_y = _q___pip_5160_1_76___block_34_tm_y;
_d___pip_5160_1_77___block_34_tm_y = _q___pip_5160_1_77___block_34_tm_y;
_d___pip_5160_1_78___block_34_tm_y = _q___pip_5160_1_78___block_34_tm_y;
_d___pip_5160_1_79___block_34_tm_y = _q___pip_5160_1_79___block_34_tm_y;
_d___pip_5160_1_80___block_34_tm_y = _q___pip_5160_1_80___block_34_tm_y;
_d___pip_5160_1_81___block_34_tm_y = _q___pip_5160_1_81___block_34_tm_y;
_d___pip_5160_1_82___block_34_tm_y = _q___pip_5160_1_82___block_34_tm_y;
_d___pip_5160_1_83___block_34_tm_y = _q___pip_5160_1_83___block_34_tm_y;
_d___pip_5160_1_84___block_34_tm_y = _q___pip_5160_1_84___block_34_tm_y;
_d___pip_5160_1_85___block_34_tm_y = _q___pip_5160_1_85___block_34_tm_y;
_d___pip_5160_1_86___block_34_tm_y = _q___pip_5160_1_86___block_34_tm_y;
_d___pip_5160_1_87___block_34_tm_y = _q___pip_5160_1_87___block_34_tm_y;
_d___pip_5160_1_88___block_34_tm_y = _q___pip_5160_1_88___block_34_tm_y;
_d___pip_5160_1_89___block_34_tm_y = _q___pip_5160_1_89___block_34_tm_y;
_d___pip_5160_1_90___block_34_tm_y = _q___pip_5160_1_90___block_34_tm_y;
_d___pip_5160_1_91___block_34_tm_y = _q___pip_5160_1_91___block_34_tm_y;
_d___pip_5160_1_92___block_34_tm_y = _q___pip_5160_1_92___block_34_tm_y;
_d___pip_5160_1_93___block_34_tm_y = _q___pip_5160_1_93___block_34_tm_y;
_d___pip_5160_1_94___block_34_tm_y = _q___pip_5160_1_94___block_34_tm_y;
_d___pip_5160_1_95___block_34_tm_y = _q___pip_5160_1_95___block_34_tm_y;
_d___pip_5160_1_96___block_34_tm_y = _q___pip_5160_1_96___block_34_tm_y;
_d___pip_5160_1_97___block_34_tm_y = _q___pip_5160_1_97___block_34_tm_y;
_d___pip_5160_1_98___block_34_tm_y = _q___pip_5160_1_98___block_34_tm_y;
_d___pip_5160_1_99___block_34_tm_y = _q___pip_5160_1_99___block_34_tm_y;
_d___pip_5160_1_100___block_34_tm_y = _q___pip_5160_1_100___block_34_tm_y;
_d___pip_5160_1_101___block_34_tm_y = _q___pip_5160_1_101___block_34_tm_y;
_d___pip_5160_1_102___block_34_tm_y = _q___pip_5160_1_102___block_34_tm_y;
_d___pip_5160_1_103___block_34_tm_y = _q___pip_5160_1_103___block_34_tm_y;
_d___pip_5160_1_104___block_34_tm_y = _q___pip_5160_1_104___block_34_tm_y;
_d___pip_5160_1_105___block_34_tm_y = _q___pip_5160_1_105___block_34_tm_y;
_d___pip_5160_1_106___block_34_tm_y = _q___pip_5160_1_106___block_34_tm_y;
_d___pip_5160_1_107___block_34_tm_y = _q___pip_5160_1_107___block_34_tm_y;
_d___pip_5160_1_108___block_34_tm_y = _q___pip_5160_1_108___block_34_tm_y;
_d___pip_5160_1_109___block_34_tm_y = _q___pip_5160_1_109___block_34_tm_y;
_d___pip_5160_1_110___block_34_tm_y = _q___pip_5160_1_110___block_34_tm_y;
_d___pip_5160_1_111___block_34_tm_y = _q___pip_5160_1_111___block_34_tm_y;
_d___pip_5160_1_112___block_34_tm_y = _q___pip_5160_1_112___block_34_tm_y;
_d___pip_5160_1_113___block_34_tm_y = _q___pip_5160_1_113___block_34_tm_y;
_d___pip_5160_1_114___block_34_tm_y = _q___pip_5160_1_114___block_34_tm_y;
_d___pip_5160_1_115___block_34_tm_y = _q___pip_5160_1_115___block_34_tm_y;
_d___pip_5160_1_116___block_34_tm_y = _q___pip_5160_1_116___block_34_tm_y;
_d___pip_5160_1_117___block_34_tm_y = _q___pip_5160_1_117___block_34_tm_y;
_d___pip_5160_1_118___block_34_tm_y = _q___pip_5160_1_118___block_34_tm_y;
_d___pip_5160_1_119___block_34_tm_y = _q___pip_5160_1_119___block_34_tm_y;
_d___pip_5160_1_120___block_34_tm_y = _q___pip_5160_1_120___block_34_tm_y;
_d___pip_5160_1_121___block_34_tm_y = _q___pip_5160_1_121___block_34_tm_y;
_d___pip_5160_1_122___block_34_tm_y = _q___pip_5160_1_122___block_34_tm_y;
_d___pip_5160_1_123___block_34_tm_y = _q___pip_5160_1_123___block_34_tm_y;
_d___pip_5160_1_124___block_34_tm_y = _q___pip_5160_1_124___block_34_tm_y;
_d___pip_5160_1_125___block_34_tm_y = _q___pip_5160_1_125___block_34_tm_y;
_d___pip_5160_1_126___block_34_tm_y = _q___pip_5160_1_126___block_34_tm_y;
_d___pip_5160_1_127___block_34_tm_y = _q___pip_5160_1_127___block_34_tm_y;
_d___pip_5160_1_128___block_34_tm_y = _q___pip_5160_1_128___block_34_tm_y;
_d___pip_5160_1_129___block_34_tm_y = _q___pip_5160_1_129___block_34_tm_y;
_d___pip_5160_1_130___block_34_tm_y = _q___pip_5160_1_130___block_34_tm_y;
_d___pip_5160_1_131___block_34_tm_y = _q___pip_5160_1_131___block_34_tm_y;
_d___pip_5160_1_132___block_34_tm_y = _q___pip_5160_1_132___block_34_tm_y;
_d___pip_5160_1_133___block_34_tm_y = _q___pip_5160_1_133___block_34_tm_y;
_d___pip_5160_1_134___block_34_tm_y = _q___pip_5160_1_134___block_34_tm_y;
_d___pip_5160_1_6___block_34_tm_z = _q___pip_5160_1_6___block_34_tm_z;
_d___pip_5160_1_7___block_34_tm_z = _q___pip_5160_1_7___block_34_tm_z;
_d___pip_5160_1_8___block_34_tm_z = _q___pip_5160_1_8___block_34_tm_z;
_d___pip_5160_1_9___block_34_tm_z = _q___pip_5160_1_9___block_34_tm_z;
_d___pip_5160_1_10___block_34_tm_z = _q___pip_5160_1_10___block_34_tm_z;
_d___pip_5160_1_11___block_34_tm_z = _q___pip_5160_1_11___block_34_tm_z;
_d___pip_5160_1_12___block_34_tm_z = _q___pip_5160_1_12___block_34_tm_z;
_d___pip_5160_1_13___block_34_tm_z = _q___pip_5160_1_13___block_34_tm_z;
_d___pip_5160_1_14___block_34_tm_z = _q___pip_5160_1_14___block_34_tm_z;
_d___pip_5160_1_15___block_34_tm_z = _q___pip_5160_1_15___block_34_tm_z;
_d___pip_5160_1_16___block_34_tm_z = _q___pip_5160_1_16___block_34_tm_z;
_d___pip_5160_1_17___block_34_tm_z = _q___pip_5160_1_17___block_34_tm_z;
_d___pip_5160_1_18___block_34_tm_z = _q___pip_5160_1_18___block_34_tm_z;
_d___pip_5160_1_19___block_34_tm_z = _q___pip_5160_1_19___block_34_tm_z;
_d___pip_5160_1_20___block_34_tm_z = _q___pip_5160_1_20___block_34_tm_z;
_d___pip_5160_1_21___block_34_tm_z = _q___pip_5160_1_21___block_34_tm_z;
_d___pip_5160_1_22___block_34_tm_z = _q___pip_5160_1_22___block_34_tm_z;
_d___pip_5160_1_23___block_34_tm_z = _q___pip_5160_1_23___block_34_tm_z;
_d___pip_5160_1_24___block_34_tm_z = _q___pip_5160_1_24___block_34_tm_z;
_d___pip_5160_1_25___block_34_tm_z = _q___pip_5160_1_25___block_34_tm_z;
_d___pip_5160_1_26___block_34_tm_z = _q___pip_5160_1_26___block_34_tm_z;
_d___pip_5160_1_27___block_34_tm_z = _q___pip_5160_1_27___block_34_tm_z;
_d___pip_5160_1_28___block_34_tm_z = _q___pip_5160_1_28___block_34_tm_z;
_d___pip_5160_1_29___block_34_tm_z = _q___pip_5160_1_29___block_34_tm_z;
_d___pip_5160_1_30___block_34_tm_z = _q___pip_5160_1_30___block_34_tm_z;
_d___pip_5160_1_31___block_34_tm_z = _q___pip_5160_1_31___block_34_tm_z;
_d___pip_5160_1_32___block_34_tm_z = _q___pip_5160_1_32___block_34_tm_z;
_d___pip_5160_1_33___block_34_tm_z = _q___pip_5160_1_33___block_34_tm_z;
_d___pip_5160_1_34___block_34_tm_z = _q___pip_5160_1_34___block_34_tm_z;
_d___pip_5160_1_35___block_34_tm_z = _q___pip_5160_1_35___block_34_tm_z;
_d___pip_5160_1_36___block_34_tm_z = _q___pip_5160_1_36___block_34_tm_z;
_d___pip_5160_1_37___block_34_tm_z = _q___pip_5160_1_37___block_34_tm_z;
_d___pip_5160_1_38___block_34_tm_z = _q___pip_5160_1_38___block_34_tm_z;
_d___pip_5160_1_39___block_34_tm_z = _q___pip_5160_1_39___block_34_tm_z;
_d___pip_5160_1_40___block_34_tm_z = _q___pip_5160_1_40___block_34_tm_z;
_d___pip_5160_1_41___block_34_tm_z = _q___pip_5160_1_41___block_34_tm_z;
_d___pip_5160_1_42___block_34_tm_z = _q___pip_5160_1_42___block_34_tm_z;
_d___pip_5160_1_43___block_34_tm_z = _q___pip_5160_1_43___block_34_tm_z;
_d___pip_5160_1_44___block_34_tm_z = _q___pip_5160_1_44___block_34_tm_z;
_d___pip_5160_1_45___block_34_tm_z = _q___pip_5160_1_45___block_34_tm_z;
_d___pip_5160_1_46___block_34_tm_z = _q___pip_5160_1_46___block_34_tm_z;
_d___pip_5160_1_47___block_34_tm_z = _q___pip_5160_1_47___block_34_tm_z;
_d___pip_5160_1_48___block_34_tm_z = _q___pip_5160_1_48___block_34_tm_z;
_d___pip_5160_1_49___block_34_tm_z = _q___pip_5160_1_49___block_34_tm_z;
_d___pip_5160_1_50___block_34_tm_z = _q___pip_5160_1_50___block_34_tm_z;
_d___pip_5160_1_51___block_34_tm_z = _q___pip_5160_1_51___block_34_tm_z;
_d___pip_5160_1_52___block_34_tm_z = _q___pip_5160_1_52___block_34_tm_z;
_d___pip_5160_1_53___block_34_tm_z = _q___pip_5160_1_53___block_34_tm_z;
_d___pip_5160_1_54___block_34_tm_z = _q___pip_5160_1_54___block_34_tm_z;
_d___pip_5160_1_55___block_34_tm_z = _q___pip_5160_1_55___block_34_tm_z;
_d___pip_5160_1_56___block_34_tm_z = _q___pip_5160_1_56___block_34_tm_z;
_d___pip_5160_1_57___block_34_tm_z = _q___pip_5160_1_57___block_34_tm_z;
_d___pip_5160_1_58___block_34_tm_z = _q___pip_5160_1_58___block_34_tm_z;
_d___pip_5160_1_59___block_34_tm_z = _q___pip_5160_1_59___block_34_tm_z;
_d___pip_5160_1_60___block_34_tm_z = _q___pip_5160_1_60___block_34_tm_z;
_d___pip_5160_1_61___block_34_tm_z = _q___pip_5160_1_61___block_34_tm_z;
_d___pip_5160_1_62___block_34_tm_z = _q___pip_5160_1_62___block_34_tm_z;
_d___pip_5160_1_63___block_34_tm_z = _q___pip_5160_1_63___block_34_tm_z;
_d___pip_5160_1_64___block_34_tm_z = _q___pip_5160_1_64___block_34_tm_z;
_d___pip_5160_1_65___block_34_tm_z = _q___pip_5160_1_65___block_34_tm_z;
_d___pip_5160_1_66___block_34_tm_z = _q___pip_5160_1_66___block_34_tm_z;
_d___pip_5160_1_67___block_34_tm_z = _q___pip_5160_1_67___block_34_tm_z;
_d___pip_5160_1_68___block_34_tm_z = _q___pip_5160_1_68___block_34_tm_z;
_d___pip_5160_1_69___block_34_tm_z = _q___pip_5160_1_69___block_34_tm_z;
_d___pip_5160_1_70___block_34_tm_z = _q___pip_5160_1_70___block_34_tm_z;
_d___pip_5160_1_71___block_34_tm_z = _q___pip_5160_1_71___block_34_tm_z;
_d___pip_5160_1_72___block_34_tm_z = _q___pip_5160_1_72___block_34_tm_z;
_d___pip_5160_1_73___block_34_tm_z = _q___pip_5160_1_73___block_34_tm_z;
_d___pip_5160_1_74___block_34_tm_z = _q___pip_5160_1_74___block_34_tm_z;
_d___pip_5160_1_75___block_34_tm_z = _q___pip_5160_1_75___block_34_tm_z;
_d___pip_5160_1_76___block_34_tm_z = _q___pip_5160_1_76___block_34_tm_z;
_d___pip_5160_1_77___block_34_tm_z = _q___pip_5160_1_77___block_34_tm_z;
_d___pip_5160_1_78___block_34_tm_z = _q___pip_5160_1_78___block_34_tm_z;
_d___pip_5160_1_79___block_34_tm_z = _q___pip_5160_1_79___block_34_tm_z;
_d___pip_5160_1_80___block_34_tm_z = _q___pip_5160_1_80___block_34_tm_z;
_d___pip_5160_1_81___block_34_tm_z = _q___pip_5160_1_81___block_34_tm_z;
_d___pip_5160_1_82___block_34_tm_z = _q___pip_5160_1_82___block_34_tm_z;
_d___pip_5160_1_83___block_34_tm_z = _q___pip_5160_1_83___block_34_tm_z;
_d___pip_5160_1_84___block_34_tm_z = _q___pip_5160_1_84___block_34_tm_z;
_d___pip_5160_1_85___block_34_tm_z = _q___pip_5160_1_85___block_34_tm_z;
_d___pip_5160_1_86___block_34_tm_z = _q___pip_5160_1_86___block_34_tm_z;
_d___pip_5160_1_87___block_34_tm_z = _q___pip_5160_1_87___block_34_tm_z;
_d___pip_5160_1_88___block_34_tm_z = _q___pip_5160_1_88___block_34_tm_z;
_d___pip_5160_1_89___block_34_tm_z = _q___pip_5160_1_89___block_34_tm_z;
_d___pip_5160_1_90___block_34_tm_z = _q___pip_5160_1_90___block_34_tm_z;
_d___pip_5160_1_91___block_34_tm_z = _q___pip_5160_1_91___block_34_tm_z;
_d___pip_5160_1_92___block_34_tm_z = _q___pip_5160_1_92___block_34_tm_z;
_d___pip_5160_1_93___block_34_tm_z = _q___pip_5160_1_93___block_34_tm_z;
_d___pip_5160_1_94___block_34_tm_z = _q___pip_5160_1_94___block_34_tm_z;
_d___pip_5160_1_95___block_34_tm_z = _q___pip_5160_1_95___block_34_tm_z;
_d___pip_5160_1_96___block_34_tm_z = _q___pip_5160_1_96___block_34_tm_z;
_d___pip_5160_1_97___block_34_tm_z = _q___pip_5160_1_97___block_34_tm_z;
_d___pip_5160_1_98___block_34_tm_z = _q___pip_5160_1_98___block_34_tm_z;
_d___pip_5160_1_99___block_34_tm_z = _q___pip_5160_1_99___block_34_tm_z;
_d___pip_5160_1_100___block_34_tm_z = _q___pip_5160_1_100___block_34_tm_z;
_d___pip_5160_1_101___block_34_tm_z = _q___pip_5160_1_101___block_34_tm_z;
_d___pip_5160_1_102___block_34_tm_z = _q___pip_5160_1_102___block_34_tm_z;
_d___pip_5160_1_103___block_34_tm_z = _q___pip_5160_1_103___block_34_tm_z;
_d___pip_5160_1_104___block_34_tm_z = _q___pip_5160_1_104___block_34_tm_z;
_d___pip_5160_1_105___block_34_tm_z = _q___pip_5160_1_105___block_34_tm_z;
_d___pip_5160_1_106___block_34_tm_z = _q___pip_5160_1_106___block_34_tm_z;
_d___pip_5160_1_107___block_34_tm_z = _q___pip_5160_1_107___block_34_tm_z;
_d___pip_5160_1_108___block_34_tm_z = _q___pip_5160_1_108___block_34_tm_z;
_d___pip_5160_1_109___block_34_tm_z = _q___pip_5160_1_109___block_34_tm_z;
_d___pip_5160_1_110___block_34_tm_z = _q___pip_5160_1_110___block_34_tm_z;
_d___pip_5160_1_111___block_34_tm_z = _q___pip_5160_1_111___block_34_tm_z;
_d___pip_5160_1_112___block_34_tm_z = _q___pip_5160_1_112___block_34_tm_z;
_d___pip_5160_1_113___block_34_tm_z = _q___pip_5160_1_113___block_34_tm_z;
_d___pip_5160_1_114___block_34_tm_z = _q___pip_5160_1_114___block_34_tm_z;
_d___pip_5160_1_115___block_34_tm_z = _q___pip_5160_1_115___block_34_tm_z;
_d___pip_5160_1_116___block_34_tm_z = _q___pip_5160_1_116___block_34_tm_z;
_d___pip_5160_1_117___block_34_tm_z = _q___pip_5160_1_117___block_34_tm_z;
_d___pip_5160_1_118___block_34_tm_z = _q___pip_5160_1_118___block_34_tm_z;
_d___pip_5160_1_119___block_34_tm_z = _q___pip_5160_1_119___block_34_tm_z;
_d___pip_5160_1_120___block_34_tm_z = _q___pip_5160_1_120___block_34_tm_z;
_d___pip_5160_1_121___block_34_tm_z = _q___pip_5160_1_121___block_34_tm_z;
_d___pip_5160_1_122___block_34_tm_z = _q___pip_5160_1_122___block_34_tm_z;
_d___pip_5160_1_123___block_34_tm_z = _q___pip_5160_1_123___block_34_tm_z;
_d___pip_5160_1_124___block_34_tm_z = _q___pip_5160_1_124___block_34_tm_z;
_d___pip_5160_1_125___block_34_tm_z = _q___pip_5160_1_125___block_34_tm_z;
_d___pip_5160_1_126___block_34_tm_z = _q___pip_5160_1_126___block_34_tm_z;
_d___pip_5160_1_127___block_34_tm_z = _q___pip_5160_1_127___block_34_tm_z;
_d___pip_5160_1_128___block_34_tm_z = _q___pip_5160_1_128___block_34_tm_z;
_d___pip_5160_1_129___block_34_tm_z = _q___pip_5160_1_129___block_34_tm_z;
_d___pip_5160_1_130___block_34_tm_z = _q___pip_5160_1_130___block_34_tm_z;
_d___pip_5160_1_131___block_34_tm_z = _q___pip_5160_1_131___block_34_tm_z;
_d___pip_5160_1_132___block_34_tm_z = _q___pip_5160_1_132___block_34_tm_z;
_d___pip_5160_1_133___block_34_tm_z = _q___pip_5160_1_133___block_34_tm_z;
_d___pip_5160_1_134___block_34_tm_z = _q___pip_5160_1_134___block_34_tm_z;
_d___pip_5160_1_6___block_40_dt_x = _q___pip_5160_1_6___block_40_dt_x;
_d___pip_5160_1_7___block_40_dt_x = _q___pip_5160_1_7___block_40_dt_x;
_d___pip_5160_1_8___block_40_dt_x = _q___pip_5160_1_8___block_40_dt_x;
_d___pip_5160_1_9___block_40_dt_x = _q___pip_5160_1_9___block_40_dt_x;
_d___pip_5160_1_10___block_40_dt_x = _q___pip_5160_1_10___block_40_dt_x;
_d___pip_5160_1_11___block_40_dt_x = _q___pip_5160_1_11___block_40_dt_x;
_d___pip_5160_1_12___block_40_dt_x = _q___pip_5160_1_12___block_40_dt_x;
_d___pip_5160_1_13___block_40_dt_x = _q___pip_5160_1_13___block_40_dt_x;
_d___pip_5160_1_14___block_40_dt_x = _q___pip_5160_1_14___block_40_dt_x;
_d___pip_5160_1_15___block_40_dt_x = _q___pip_5160_1_15___block_40_dt_x;
_d___pip_5160_1_16___block_40_dt_x = _q___pip_5160_1_16___block_40_dt_x;
_d___pip_5160_1_17___block_40_dt_x = _q___pip_5160_1_17___block_40_dt_x;
_d___pip_5160_1_18___block_40_dt_x = _q___pip_5160_1_18___block_40_dt_x;
_d___pip_5160_1_19___block_40_dt_x = _q___pip_5160_1_19___block_40_dt_x;
_d___pip_5160_1_20___block_40_dt_x = _q___pip_5160_1_20___block_40_dt_x;
_d___pip_5160_1_21___block_40_dt_x = _q___pip_5160_1_21___block_40_dt_x;
_d___pip_5160_1_22___block_40_dt_x = _q___pip_5160_1_22___block_40_dt_x;
_d___pip_5160_1_23___block_40_dt_x = _q___pip_5160_1_23___block_40_dt_x;
_d___pip_5160_1_24___block_40_dt_x = _q___pip_5160_1_24___block_40_dt_x;
_d___pip_5160_1_25___block_40_dt_x = _q___pip_5160_1_25___block_40_dt_x;
_d___pip_5160_1_26___block_40_dt_x = _q___pip_5160_1_26___block_40_dt_x;
_d___pip_5160_1_27___block_40_dt_x = _q___pip_5160_1_27___block_40_dt_x;
_d___pip_5160_1_28___block_40_dt_x = _q___pip_5160_1_28___block_40_dt_x;
_d___pip_5160_1_29___block_40_dt_x = _q___pip_5160_1_29___block_40_dt_x;
_d___pip_5160_1_30___block_40_dt_x = _q___pip_5160_1_30___block_40_dt_x;
_d___pip_5160_1_31___block_40_dt_x = _q___pip_5160_1_31___block_40_dt_x;
_d___pip_5160_1_32___block_40_dt_x = _q___pip_5160_1_32___block_40_dt_x;
_d___pip_5160_1_33___block_40_dt_x = _q___pip_5160_1_33___block_40_dt_x;
_d___pip_5160_1_34___block_40_dt_x = _q___pip_5160_1_34___block_40_dt_x;
_d___pip_5160_1_35___block_40_dt_x = _q___pip_5160_1_35___block_40_dt_x;
_d___pip_5160_1_36___block_40_dt_x = _q___pip_5160_1_36___block_40_dt_x;
_d___pip_5160_1_37___block_40_dt_x = _q___pip_5160_1_37___block_40_dt_x;
_d___pip_5160_1_38___block_40_dt_x = _q___pip_5160_1_38___block_40_dt_x;
_d___pip_5160_1_39___block_40_dt_x = _q___pip_5160_1_39___block_40_dt_x;
_d___pip_5160_1_40___block_40_dt_x = _q___pip_5160_1_40___block_40_dt_x;
_d___pip_5160_1_41___block_40_dt_x = _q___pip_5160_1_41___block_40_dt_x;
_d___pip_5160_1_42___block_40_dt_x = _q___pip_5160_1_42___block_40_dt_x;
_d___pip_5160_1_43___block_40_dt_x = _q___pip_5160_1_43___block_40_dt_x;
_d___pip_5160_1_44___block_40_dt_x = _q___pip_5160_1_44___block_40_dt_x;
_d___pip_5160_1_45___block_40_dt_x = _q___pip_5160_1_45___block_40_dt_x;
_d___pip_5160_1_46___block_40_dt_x = _q___pip_5160_1_46___block_40_dt_x;
_d___pip_5160_1_47___block_40_dt_x = _q___pip_5160_1_47___block_40_dt_x;
_d___pip_5160_1_48___block_40_dt_x = _q___pip_5160_1_48___block_40_dt_x;
_d___pip_5160_1_49___block_40_dt_x = _q___pip_5160_1_49___block_40_dt_x;
_d___pip_5160_1_50___block_40_dt_x = _q___pip_5160_1_50___block_40_dt_x;
_d___pip_5160_1_51___block_40_dt_x = _q___pip_5160_1_51___block_40_dt_x;
_d___pip_5160_1_52___block_40_dt_x = _q___pip_5160_1_52___block_40_dt_x;
_d___pip_5160_1_53___block_40_dt_x = _q___pip_5160_1_53___block_40_dt_x;
_d___pip_5160_1_54___block_40_dt_x = _q___pip_5160_1_54___block_40_dt_x;
_d___pip_5160_1_55___block_40_dt_x = _q___pip_5160_1_55___block_40_dt_x;
_d___pip_5160_1_56___block_40_dt_x = _q___pip_5160_1_56___block_40_dt_x;
_d___pip_5160_1_57___block_40_dt_x = _q___pip_5160_1_57___block_40_dt_x;
_d___pip_5160_1_58___block_40_dt_x = _q___pip_5160_1_58___block_40_dt_x;
_d___pip_5160_1_59___block_40_dt_x = _q___pip_5160_1_59___block_40_dt_x;
_d___pip_5160_1_60___block_40_dt_x = _q___pip_5160_1_60___block_40_dt_x;
_d___pip_5160_1_61___block_40_dt_x = _q___pip_5160_1_61___block_40_dt_x;
_d___pip_5160_1_62___block_40_dt_x = _q___pip_5160_1_62___block_40_dt_x;
_d___pip_5160_1_63___block_40_dt_x = _q___pip_5160_1_63___block_40_dt_x;
_d___pip_5160_1_64___block_40_dt_x = _q___pip_5160_1_64___block_40_dt_x;
_d___pip_5160_1_65___block_40_dt_x = _q___pip_5160_1_65___block_40_dt_x;
_d___pip_5160_1_66___block_40_dt_x = _q___pip_5160_1_66___block_40_dt_x;
_d___pip_5160_1_67___block_40_dt_x = _q___pip_5160_1_67___block_40_dt_x;
_d___pip_5160_1_68___block_40_dt_x = _q___pip_5160_1_68___block_40_dt_x;
_d___pip_5160_1_69___block_40_dt_x = _q___pip_5160_1_69___block_40_dt_x;
_d___pip_5160_1_70___block_40_dt_x = _q___pip_5160_1_70___block_40_dt_x;
_d___pip_5160_1_71___block_40_dt_x = _q___pip_5160_1_71___block_40_dt_x;
_d___pip_5160_1_72___block_40_dt_x = _q___pip_5160_1_72___block_40_dt_x;
_d___pip_5160_1_73___block_40_dt_x = _q___pip_5160_1_73___block_40_dt_x;
_d___pip_5160_1_74___block_40_dt_x = _q___pip_5160_1_74___block_40_dt_x;
_d___pip_5160_1_75___block_40_dt_x = _q___pip_5160_1_75___block_40_dt_x;
_d___pip_5160_1_76___block_40_dt_x = _q___pip_5160_1_76___block_40_dt_x;
_d___pip_5160_1_77___block_40_dt_x = _q___pip_5160_1_77___block_40_dt_x;
_d___pip_5160_1_78___block_40_dt_x = _q___pip_5160_1_78___block_40_dt_x;
_d___pip_5160_1_79___block_40_dt_x = _q___pip_5160_1_79___block_40_dt_x;
_d___pip_5160_1_80___block_40_dt_x = _q___pip_5160_1_80___block_40_dt_x;
_d___pip_5160_1_81___block_40_dt_x = _q___pip_5160_1_81___block_40_dt_x;
_d___pip_5160_1_82___block_40_dt_x = _q___pip_5160_1_82___block_40_dt_x;
_d___pip_5160_1_83___block_40_dt_x = _q___pip_5160_1_83___block_40_dt_x;
_d___pip_5160_1_84___block_40_dt_x = _q___pip_5160_1_84___block_40_dt_x;
_d___pip_5160_1_85___block_40_dt_x = _q___pip_5160_1_85___block_40_dt_x;
_d___pip_5160_1_86___block_40_dt_x = _q___pip_5160_1_86___block_40_dt_x;
_d___pip_5160_1_87___block_40_dt_x = _q___pip_5160_1_87___block_40_dt_x;
_d___pip_5160_1_88___block_40_dt_x = _q___pip_5160_1_88___block_40_dt_x;
_d___pip_5160_1_89___block_40_dt_x = _q___pip_5160_1_89___block_40_dt_x;
_d___pip_5160_1_90___block_40_dt_x = _q___pip_5160_1_90___block_40_dt_x;
_d___pip_5160_1_91___block_40_dt_x = _q___pip_5160_1_91___block_40_dt_x;
_d___pip_5160_1_92___block_40_dt_x = _q___pip_5160_1_92___block_40_dt_x;
_d___pip_5160_1_93___block_40_dt_x = _q___pip_5160_1_93___block_40_dt_x;
_d___pip_5160_1_94___block_40_dt_x = _q___pip_5160_1_94___block_40_dt_x;
_d___pip_5160_1_95___block_40_dt_x = _q___pip_5160_1_95___block_40_dt_x;
_d___pip_5160_1_96___block_40_dt_x = _q___pip_5160_1_96___block_40_dt_x;
_d___pip_5160_1_97___block_40_dt_x = _q___pip_5160_1_97___block_40_dt_x;
_d___pip_5160_1_98___block_40_dt_x = _q___pip_5160_1_98___block_40_dt_x;
_d___pip_5160_1_99___block_40_dt_x = _q___pip_5160_1_99___block_40_dt_x;
_d___pip_5160_1_100___block_40_dt_x = _q___pip_5160_1_100___block_40_dt_x;
_d___pip_5160_1_101___block_40_dt_x = _q___pip_5160_1_101___block_40_dt_x;
_d___pip_5160_1_102___block_40_dt_x = _q___pip_5160_1_102___block_40_dt_x;
_d___pip_5160_1_103___block_40_dt_x = _q___pip_5160_1_103___block_40_dt_x;
_d___pip_5160_1_104___block_40_dt_x = _q___pip_5160_1_104___block_40_dt_x;
_d___pip_5160_1_105___block_40_dt_x = _q___pip_5160_1_105___block_40_dt_x;
_d___pip_5160_1_106___block_40_dt_x = _q___pip_5160_1_106___block_40_dt_x;
_d___pip_5160_1_107___block_40_dt_x = _q___pip_5160_1_107___block_40_dt_x;
_d___pip_5160_1_108___block_40_dt_x = _q___pip_5160_1_108___block_40_dt_x;
_d___pip_5160_1_109___block_40_dt_x = _q___pip_5160_1_109___block_40_dt_x;
_d___pip_5160_1_110___block_40_dt_x = _q___pip_5160_1_110___block_40_dt_x;
_d___pip_5160_1_111___block_40_dt_x = _q___pip_5160_1_111___block_40_dt_x;
_d___pip_5160_1_112___block_40_dt_x = _q___pip_5160_1_112___block_40_dt_x;
_d___pip_5160_1_113___block_40_dt_x = _q___pip_5160_1_113___block_40_dt_x;
_d___pip_5160_1_114___block_40_dt_x = _q___pip_5160_1_114___block_40_dt_x;
_d___pip_5160_1_115___block_40_dt_x = _q___pip_5160_1_115___block_40_dt_x;
_d___pip_5160_1_116___block_40_dt_x = _q___pip_5160_1_116___block_40_dt_x;
_d___pip_5160_1_117___block_40_dt_x = _q___pip_5160_1_117___block_40_dt_x;
_d___pip_5160_1_118___block_40_dt_x = _q___pip_5160_1_118___block_40_dt_x;
_d___pip_5160_1_119___block_40_dt_x = _q___pip_5160_1_119___block_40_dt_x;
_d___pip_5160_1_120___block_40_dt_x = _q___pip_5160_1_120___block_40_dt_x;
_d___pip_5160_1_121___block_40_dt_x = _q___pip_5160_1_121___block_40_dt_x;
_d___pip_5160_1_122___block_40_dt_x = _q___pip_5160_1_122___block_40_dt_x;
_d___pip_5160_1_123___block_40_dt_x = _q___pip_5160_1_123___block_40_dt_x;
_d___pip_5160_1_124___block_40_dt_x = _q___pip_5160_1_124___block_40_dt_x;
_d___pip_5160_1_125___block_40_dt_x = _q___pip_5160_1_125___block_40_dt_x;
_d___pip_5160_1_126___block_40_dt_x = _q___pip_5160_1_126___block_40_dt_x;
_d___pip_5160_1_127___block_40_dt_x = _q___pip_5160_1_127___block_40_dt_x;
_d___pip_5160_1_128___block_40_dt_x = _q___pip_5160_1_128___block_40_dt_x;
_d___pip_5160_1_129___block_40_dt_x = _q___pip_5160_1_129___block_40_dt_x;
_d___pip_5160_1_130___block_40_dt_x = _q___pip_5160_1_130___block_40_dt_x;
_d___pip_5160_1_131___block_40_dt_x = _q___pip_5160_1_131___block_40_dt_x;
_d___pip_5160_1_132___block_40_dt_x = _q___pip_5160_1_132___block_40_dt_x;
_d___pip_5160_1_133___block_40_dt_x = _q___pip_5160_1_133___block_40_dt_x;
_d___pip_5160_1_134___block_40_dt_x = _q___pip_5160_1_134___block_40_dt_x;
_d___pip_5160_1_6___block_40_dt_y = _q___pip_5160_1_6___block_40_dt_y;
_d___pip_5160_1_7___block_40_dt_y = _q___pip_5160_1_7___block_40_dt_y;
_d___pip_5160_1_8___block_40_dt_y = _q___pip_5160_1_8___block_40_dt_y;
_d___pip_5160_1_9___block_40_dt_y = _q___pip_5160_1_9___block_40_dt_y;
_d___pip_5160_1_10___block_40_dt_y = _q___pip_5160_1_10___block_40_dt_y;
_d___pip_5160_1_11___block_40_dt_y = _q___pip_5160_1_11___block_40_dt_y;
_d___pip_5160_1_12___block_40_dt_y = _q___pip_5160_1_12___block_40_dt_y;
_d___pip_5160_1_13___block_40_dt_y = _q___pip_5160_1_13___block_40_dt_y;
_d___pip_5160_1_14___block_40_dt_y = _q___pip_5160_1_14___block_40_dt_y;
_d___pip_5160_1_15___block_40_dt_y = _q___pip_5160_1_15___block_40_dt_y;
_d___pip_5160_1_16___block_40_dt_y = _q___pip_5160_1_16___block_40_dt_y;
_d___pip_5160_1_17___block_40_dt_y = _q___pip_5160_1_17___block_40_dt_y;
_d___pip_5160_1_18___block_40_dt_y = _q___pip_5160_1_18___block_40_dt_y;
_d___pip_5160_1_19___block_40_dt_y = _q___pip_5160_1_19___block_40_dt_y;
_d___pip_5160_1_20___block_40_dt_y = _q___pip_5160_1_20___block_40_dt_y;
_d___pip_5160_1_21___block_40_dt_y = _q___pip_5160_1_21___block_40_dt_y;
_d___pip_5160_1_22___block_40_dt_y = _q___pip_5160_1_22___block_40_dt_y;
_d___pip_5160_1_23___block_40_dt_y = _q___pip_5160_1_23___block_40_dt_y;
_d___pip_5160_1_24___block_40_dt_y = _q___pip_5160_1_24___block_40_dt_y;
_d___pip_5160_1_25___block_40_dt_y = _q___pip_5160_1_25___block_40_dt_y;
_d___pip_5160_1_26___block_40_dt_y = _q___pip_5160_1_26___block_40_dt_y;
_d___pip_5160_1_27___block_40_dt_y = _q___pip_5160_1_27___block_40_dt_y;
_d___pip_5160_1_28___block_40_dt_y = _q___pip_5160_1_28___block_40_dt_y;
_d___pip_5160_1_29___block_40_dt_y = _q___pip_5160_1_29___block_40_dt_y;
_d___pip_5160_1_30___block_40_dt_y = _q___pip_5160_1_30___block_40_dt_y;
_d___pip_5160_1_31___block_40_dt_y = _q___pip_5160_1_31___block_40_dt_y;
_d___pip_5160_1_32___block_40_dt_y = _q___pip_5160_1_32___block_40_dt_y;
_d___pip_5160_1_33___block_40_dt_y = _q___pip_5160_1_33___block_40_dt_y;
_d___pip_5160_1_34___block_40_dt_y = _q___pip_5160_1_34___block_40_dt_y;
_d___pip_5160_1_35___block_40_dt_y = _q___pip_5160_1_35___block_40_dt_y;
_d___pip_5160_1_36___block_40_dt_y = _q___pip_5160_1_36___block_40_dt_y;
_d___pip_5160_1_37___block_40_dt_y = _q___pip_5160_1_37___block_40_dt_y;
_d___pip_5160_1_38___block_40_dt_y = _q___pip_5160_1_38___block_40_dt_y;
_d___pip_5160_1_39___block_40_dt_y = _q___pip_5160_1_39___block_40_dt_y;
_d___pip_5160_1_40___block_40_dt_y = _q___pip_5160_1_40___block_40_dt_y;
_d___pip_5160_1_41___block_40_dt_y = _q___pip_5160_1_41___block_40_dt_y;
_d___pip_5160_1_42___block_40_dt_y = _q___pip_5160_1_42___block_40_dt_y;
_d___pip_5160_1_43___block_40_dt_y = _q___pip_5160_1_43___block_40_dt_y;
_d___pip_5160_1_44___block_40_dt_y = _q___pip_5160_1_44___block_40_dt_y;
_d___pip_5160_1_45___block_40_dt_y = _q___pip_5160_1_45___block_40_dt_y;
_d___pip_5160_1_46___block_40_dt_y = _q___pip_5160_1_46___block_40_dt_y;
_d___pip_5160_1_47___block_40_dt_y = _q___pip_5160_1_47___block_40_dt_y;
_d___pip_5160_1_48___block_40_dt_y = _q___pip_5160_1_48___block_40_dt_y;
_d___pip_5160_1_49___block_40_dt_y = _q___pip_5160_1_49___block_40_dt_y;
_d___pip_5160_1_50___block_40_dt_y = _q___pip_5160_1_50___block_40_dt_y;
_d___pip_5160_1_51___block_40_dt_y = _q___pip_5160_1_51___block_40_dt_y;
_d___pip_5160_1_52___block_40_dt_y = _q___pip_5160_1_52___block_40_dt_y;
_d___pip_5160_1_53___block_40_dt_y = _q___pip_5160_1_53___block_40_dt_y;
_d___pip_5160_1_54___block_40_dt_y = _q___pip_5160_1_54___block_40_dt_y;
_d___pip_5160_1_55___block_40_dt_y = _q___pip_5160_1_55___block_40_dt_y;
_d___pip_5160_1_56___block_40_dt_y = _q___pip_5160_1_56___block_40_dt_y;
_d___pip_5160_1_57___block_40_dt_y = _q___pip_5160_1_57___block_40_dt_y;
_d___pip_5160_1_58___block_40_dt_y = _q___pip_5160_1_58___block_40_dt_y;
_d___pip_5160_1_59___block_40_dt_y = _q___pip_5160_1_59___block_40_dt_y;
_d___pip_5160_1_60___block_40_dt_y = _q___pip_5160_1_60___block_40_dt_y;
_d___pip_5160_1_61___block_40_dt_y = _q___pip_5160_1_61___block_40_dt_y;
_d___pip_5160_1_62___block_40_dt_y = _q___pip_5160_1_62___block_40_dt_y;
_d___pip_5160_1_63___block_40_dt_y = _q___pip_5160_1_63___block_40_dt_y;
_d___pip_5160_1_64___block_40_dt_y = _q___pip_5160_1_64___block_40_dt_y;
_d___pip_5160_1_65___block_40_dt_y = _q___pip_5160_1_65___block_40_dt_y;
_d___pip_5160_1_66___block_40_dt_y = _q___pip_5160_1_66___block_40_dt_y;
_d___pip_5160_1_67___block_40_dt_y = _q___pip_5160_1_67___block_40_dt_y;
_d___pip_5160_1_68___block_40_dt_y = _q___pip_5160_1_68___block_40_dt_y;
_d___pip_5160_1_69___block_40_dt_y = _q___pip_5160_1_69___block_40_dt_y;
_d___pip_5160_1_70___block_40_dt_y = _q___pip_5160_1_70___block_40_dt_y;
_d___pip_5160_1_71___block_40_dt_y = _q___pip_5160_1_71___block_40_dt_y;
_d___pip_5160_1_72___block_40_dt_y = _q___pip_5160_1_72___block_40_dt_y;
_d___pip_5160_1_73___block_40_dt_y = _q___pip_5160_1_73___block_40_dt_y;
_d___pip_5160_1_74___block_40_dt_y = _q___pip_5160_1_74___block_40_dt_y;
_d___pip_5160_1_75___block_40_dt_y = _q___pip_5160_1_75___block_40_dt_y;
_d___pip_5160_1_76___block_40_dt_y = _q___pip_5160_1_76___block_40_dt_y;
_d___pip_5160_1_77___block_40_dt_y = _q___pip_5160_1_77___block_40_dt_y;
_d___pip_5160_1_78___block_40_dt_y = _q___pip_5160_1_78___block_40_dt_y;
_d___pip_5160_1_79___block_40_dt_y = _q___pip_5160_1_79___block_40_dt_y;
_d___pip_5160_1_80___block_40_dt_y = _q___pip_5160_1_80___block_40_dt_y;
_d___pip_5160_1_81___block_40_dt_y = _q___pip_5160_1_81___block_40_dt_y;
_d___pip_5160_1_82___block_40_dt_y = _q___pip_5160_1_82___block_40_dt_y;
_d___pip_5160_1_83___block_40_dt_y = _q___pip_5160_1_83___block_40_dt_y;
_d___pip_5160_1_84___block_40_dt_y = _q___pip_5160_1_84___block_40_dt_y;
_d___pip_5160_1_85___block_40_dt_y = _q___pip_5160_1_85___block_40_dt_y;
_d___pip_5160_1_86___block_40_dt_y = _q___pip_5160_1_86___block_40_dt_y;
_d___pip_5160_1_87___block_40_dt_y = _q___pip_5160_1_87___block_40_dt_y;
_d___pip_5160_1_88___block_40_dt_y = _q___pip_5160_1_88___block_40_dt_y;
_d___pip_5160_1_89___block_40_dt_y = _q___pip_5160_1_89___block_40_dt_y;
_d___pip_5160_1_90___block_40_dt_y = _q___pip_5160_1_90___block_40_dt_y;
_d___pip_5160_1_91___block_40_dt_y = _q___pip_5160_1_91___block_40_dt_y;
_d___pip_5160_1_92___block_40_dt_y = _q___pip_5160_1_92___block_40_dt_y;
_d___pip_5160_1_93___block_40_dt_y = _q___pip_5160_1_93___block_40_dt_y;
_d___pip_5160_1_94___block_40_dt_y = _q___pip_5160_1_94___block_40_dt_y;
_d___pip_5160_1_95___block_40_dt_y = _q___pip_5160_1_95___block_40_dt_y;
_d___pip_5160_1_96___block_40_dt_y = _q___pip_5160_1_96___block_40_dt_y;
_d___pip_5160_1_97___block_40_dt_y = _q___pip_5160_1_97___block_40_dt_y;
_d___pip_5160_1_98___block_40_dt_y = _q___pip_5160_1_98___block_40_dt_y;
_d___pip_5160_1_99___block_40_dt_y = _q___pip_5160_1_99___block_40_dt_y;
_d___pip_5160_1_100___block_40_dt_y = _q___pip_5160_1_100___block_40_dt_y;
_d___pip_5160_1_101___block_40_dt_y = _q___pip_5160_1_101___block_40_dt_y;
_d___pip_5160_1_102___block_40_dt_y = _q___pip_5160_1_102___block_40_dt_y;
_d___pip_5160_1_103___block_40_dt_y = _q___pip_5160_1_103___block_40_dt_y;
_d___pip_5160_1_104___block_40_dt_y = _q___pip_5160_1_104___block_40_dt_y;
_d___pip_5160_1_105___block_40_dt_y = _q___pip_5160_1_105___block_40_dt_y;
_d___pip_5160_1_106___block_40_dt_y = _q___pip_5160_1_106___block_40_dt_y;
_d___pip_5160_1_107___block_40_dt_y = _q___pip_5160_1_107___block_40_dt_y;
_d___pip_5160_1_108___block_40_dt_y = _q___pip_5160_1_108___block_40_dt_y;
_d___pip_5160_1_109___block_40_dt_y = _q___pip_5160_1_109___block_40_dt_y;
_d___pip_5160_1_110___block_40_dt_y = _q___pip_5160_1_110___block_40_dt_y;
_d___pip_5160_1_111___block_40_dt_y = _q___pip_5160_1_111___block_40_dt_y;
_d___pip_5160_1_112___block_40_dt_y = _q___pip_5160_1_112___block_40_dt_y;
_d___pip_5160_1_113___block_40_dt_y = _q___pip_5160_1_113___block_40_dt_y;
_d___pip_5160_1_114___block_40_dt_y = _q___pip_5160_1_114___block_40_dt_y;
_d___pip_5160_1_115___block_40_dt_y = _q___pip_5160_1_115___block_40_dt_y;
_d___pip_5160_1_116___block_40_dt_y = _q___pip_5160_1_116___block_40_dt_y;
_d___pip_5160_1_117___block_40_dt_y = _q___pip_5160_1_117___block_40_dt_y;
_d___pip_5160_1_118___block_40_dt_y = _q___pip_5160_1_118___block_40_dt_y;
_d___pip_5160_1_119___block_40_dt_y = _q___pip_5160_1_119___block_40_dt_y;
_d___pip_5160_1_120___block_40_dt_y = _q___pip_5160_1_120___block_40_dt_y;
_d___pip_5160_1_121___block_40_dt_y = _q___pip_5160_1_121___block_40_dt_y;
_d___pip_5160_1_122___block_40_dt_y = _q___pip_5160_1_122___block_40_dt_y;
_d___pip_5160_1_123___block_40_dt_y = _q___pip_5160_1_123___block_40_dt_y;
_d___pip_5160_1_124___block_40_dt_y = _q___pip_5160_1_124___block_40_dt_y;
_d___pip_5160_1_125___block_40_dt_y = _q___pip_5160_1_125___block_40_dt_y;
_d___pip_5160_1_126___block_40_dt_y = _q___pip_5160_1_126___block_40_dt_y;
_d___pip_5160_1_127___block_40_dt_y = _q___pip_5160_1_127___block_40_dt_y;
_d___pip_5160_1_128___block_40_dt_y = _q___pip_5160_1_128___block_40_dt_y;
_d___pip_5160_1_129___block_40_dt_y = _q___pip_5160_1_129___block_40_dt_y;
_d___pip_5160_1_130___block_40_dt_y = _q___pip_5160_1_130___block_40_dt_y;
_d___pip_5160_1_131___block_40_dt_y = _q___pip_5160_1_131___block_40_dt_y;
_d___pip_5160_1_132___block_40_dt_y = _q___pip_5160_1_132___block_40_dt_y;
_d___pip_5160_1_133___block_40_dt_y = _q___pip_5160_1_133___block_40_dt_y;
_d___pip_5160_1_134___block_40_dt_y = _q___pip_5160_1_134___block_40_dt_y;
_d___pip_5160_1_6___block_40_dt_z = _q___pip_5160_1_6___block_40_dt_z;
_d___pip_5160_1_7___block_40_dt_z = _q___pip_5160_1_7___block_40_dt_z;
_d___pip_5160_1_8___block_40_dt_z = _q___pip_5160_1_8___block_40_dt_z;
_d___pip_5160_1_9___block_40_dt_z = _q___pip_5160_1_9___block_40_dt_z;
_d___pip_5160_1_10___block_40_dt_z = _q___pip_5160_1_10___block_40_dt_z;
_d___pip_5160_1_11___block_40_dt_z = _q___pip_5160_1_11___block_40_dt_z;
_d___pip_5160_1_12___block_40_dt_z = _q___pip_5160_1_12___block_40_dt_z;
_d___pip_5160_1_13___block_40_dt_z = _q___pip_5160_1_13___block_40_dt_z;
_d___pip_5160_1_14___block_40_dt_z = _q___pip_5160_1_14___block_40_dt_z;
_d___pip_5160_1_15___block_40_dt_z = _q___pip_5160_1_15___block_40_dt_z;
_d___pip_5160_1_16___block_40_dt_z = _q___pip_5160_1_16___block_40_dt_z;
_d___pip_5160_1_17___block_40_dt_z = _q___pip_5160_1_17___block_40_dt_z;
_d___pip_5160_1_18___block_40_dt_z = _q___pip_5160_1_18___block_40_dt_z;
_d___pip_5160_1_19___block_40_dt_z = _q___pip_5160_1_19___block_40_dt_z;
_d___pip_5160_1_20___block_40_dt_z = _q___pip_5160_1_20___block_40_dt_z;
_d___pip_5160_1_21___block_40_dt_z = _q___pip_5160_1_21___block_40_dt_z;
_d___pip_5160_1_22___block_40_dt_z = _q___pip_5160_1_22___block_40_dt_z;
_d___pip_5160_1_23___block_40_dt_z = _q___pip_5160_1_23___block_40_dt_z;
_d___pip_5160_1_24___block_40_dt_z = _q___pip_5160_1_24___block_40_dt_z;
_d___pip_5160_1_25___block_40_dt_z = _q___pip_5160_1_25___block_40_dt_z;
_d___pip_5160_1_26___block_40_dt_z = _q___pip_5160_1_26___block_40_dt_z;
_d___pip_5160_1_27___block_40_dt_z = _q___pip_5160_1_27___block_40_dt_z;
_d___pip_5160_1_28___block_40_dt_z = _q___pip_5160_1_28___block_40_dt_z;
_d___pip_5160_1_29___block_40_dt_z = _q___pip_5160_1_29___block_40_dt_z;
_d___pip_5160_1_30___block_40_dt_z = _q___pip_5160_1_30___block_40_dt_z;
_d___pip_5160_1_31___block_40_dt_z = _q___pip_5160_1_31___block_40_dt_z;
_d___pip_5160_1_32___block_40_dt_z = _q___pip_5160_1_32___block_40_dt_z;
_d___pip_5160_1_33___block_40_dt_z = _q___pip_5160_1_33___block_40_dt_z;
_d___pip_5160_1_34___block_40_dt_z = _q___pip_5160_1_34___block_40_dt_z;
_d___pip_5160_1_35___block_40_dt_z = _q___pip_5160_1_35___block_40_dt_z;
_d___pip_5160_1_36___block_40_dt_z = _q___pip_5160_1_36___block_40_dt_z;
_d___pip_5160_1_37___block_40_dt_z = _q___pip_5160_1_37___block_40_dt_z;
_d___pip_5160_1_38___block_40_dt_z = _q___pip_5160_1_38___block_40_dt_z;
_d___pip_5160_1_39___block_40_dt_z = _q___pip_5160_1_39___block_40_dt_z;
_d___pip_5160_1_40___block_40_dt_z = _q___pip_5160_1_40___block_40_dt_z;
_d___pip_5160_1_41___block_40_dt_z = _q___pip_5160_1_41___block_40_dt_z;
_d___pip_5160_1_42___block_40_dt_z = _q___pip_5160_1_42___block_40_dt_z;
_d___pip_5160_1_43___block_40_dt_z = _q___pip_5160_1_43___block_40_dt_z;
_d___pip_5160_1_44___block_40_dt_z = _q___pip_5160_1_44___block_40_dt_z;
_d___pip_5160_1_45___block_40_dt_z = _q___pip_5160_1_45___block_40_dt_z;
_d___pip_5160_1_46___block_40_dt_z = _q___pip_5160_1_46___block_40_dt_z;
_d___pip_5160_1_47___block_40_dt_z = _q___pip_5160_1_47___block_40_dt_z;
_d___pip_5160_1_48___block_40_dt_z = _q___pip_5160_1_48___block_40_dt_z;
_d___pip_5160_1_49___block_40_dt_z = _q___pip_5160_1_49___block_40_dt_z;
_d___pip_5160_1_50___block_40_dt_z = _q___pip_5160_1_50___block_40_dt_z;
_d___pip_5160_1_51___block_40_dt_z = _q___pip_5160_1_51___block_40_dt_z;
_d___pip_5160_1_52___block_40_dt_z = _q___pip_5160_1_52___block_40_dt_z;
_d___pip_5160_1_53___block_40_dt_z = _q___pip_5160_1_53___block_40_dt_z;
_d___pip_5160_1_54___block_40_dt_z = _q___pip_5160_1_54___block_40_dt_z;
_d___pip_5160_1_55___block_40_dt_z = _q___pip_5160_1_55___block_40_dt_z;
_d___pip_5160_1_56___block_40_dt_z = _q___pip_5160_1_56___block_40_dt_z;
_d___pip_5160_1_57___block_40_dt_z = _q___pip_5160_1_57___block_40_dt_z;
_d___pip_5160_1_58___block_40_dt_z = _q___pip_5160_1_58___block_40_dt_z;
_d___pip_5160_1_59___block_40_dt_z = _q___pip_5160_1_59___block_40_dt_z;
_d___pip_5160_1_60___block_40_dt_z = _q___pip_5160_1_60___block_40_dt_z;
_d___pip_5160_1_61___block_40_dt_z = _q___pip_5160_1_61___block_40_dt_z;
_d___pip_5160_1_62___block_40_dt_z = _q___pip_5160_1_62___block_40_dt_z;
_d___pip_5160_1_63___block_40_dt_z = _q___pip_5160_1_63___block_40_dt_z;
_d___pip_5160_1_64___block_40_dt_z = _q___pip_5160_1_64___block_40_dt_z;
_d___pip_5160_1_65___block_40_dt_z = _q___pip_5160_1_65___block_40_dt_z;
_d___pip_5160_1_66___block_40_dt_z = _q___pip_5160_1_66___block_40_dt_z;
_d___pip_5160_1_67___block_40_dt_z = _q___pip_5160_1_67___block_40_dt_z;
_d___pip_5160_1_68___block_40_dt_z = _q___pip_5160_1_68___block_40_dt_z;
_d___pip_5160_1_69___block_40_dt_z = _q___pip_5160_1_69___block_40_dt_z;
_d___pip_5160_1_70___block_40_dt_z = _q___pip_5160_1_70___block_40_dt_z;
_d___pip_5160_1_71___block_40_dt_z = _q___pip_5160_1_71___block_40_dt_z;
_d___pip_5160_1_72___block_40_dt_z = _q___pip_5160_1_72___block_40_dt_z;
_d___pip_5160_1_73___block_40_dt_z = _q___pip_5160_1_73___block_40_dt_z;
_d___pip_5160_1_74___block_40_dt_z = _q___pip_5160_1_74___block_40_dt_z;
_d___pip_5160_1_75___block_40_dt_z = _q___pip_5160_1_75___block_40_dt_z;
_d___pip_5160_1_76___block_40_dt_z = _q___pip_5160_1_76___block_40_dt_z;
_d___pip_5160_1_77___block_40_dt_z = _q___pip_5160_1_77___block_40_dt_z;
_d___pip_5160_1_78___block_40_dt_z = _q___pip_5160_1_78___block_40_dt_z;
_d___pip_5160_1_79___block_40_dt_z = _q___pip_5160_1_79___block_40_dt_z;
_d___pip_5160_1_80___block_40_dt_z = _q___pip_5160_1_80___block_40_dt_z;
_d___pip_5160_1_81___block_40_dt_z = _q___pip_5160_1_81___block_40_dt_z;
_d___pip_5160_1_82___block_40_dt_z = _q___pip_5160_1_82___block_40_dt_z;
_d___pip_5160_1_83___block_40_dt_z = _q___pip_5160_1_83___block_40_dt_z;
_d___pip_5160_1_84___block_40_dt_z = _q___pip_5160_1_84___block_40_dt_z;
_d___pip_5160_1_85___block_40_dt_z = _q___pip_5160_1_85___block_40_dt_z;
_d___pip_5160_1_86___block_40_dt_z = _q___pip_5160_1_86___block_40_dt_z;
_d___pip_5160_1_87___block_40_dt_z = _q___pip_5160_1_87___block_40_dt_z;
_d___pip_5160_1_88___block_40_dt_z = _q___pip_5160_1_88___block_40_dt_z;
_d___pip_5160_1_89___block_40_dt_z = _q___pip_5160_1_89___block_40_dt_z;
_d___pip_5160_1_90___block_40_dt_z = _q___pip_5160_1_90___block_40_dt_z;
_d___pip_5160_1_91___block_40_dt_z = _q___pip_5160_1_91___block_40_dt_z;
_d___pip_5160_1_92___block_40_dt_z = _q___pip_5160_1_92___block_40_dt_z;
_d___pip_5160_1_93___block_40_dt_z = _q___pip_5160_1_93___block_40_dt_z;
_d___pip_5160_1_94___block_40_dt_z = _q___pip_5160_1_94___block_40_dt_z;
_d___pip_5160_1_95___block_40_dt_z = _q___pip_5160_1_95___block_40_dt_z;
_d___pip_5160_1_96___block_40_dt_z = _q___pip_5160_1_96___block_40_dt_z;
_d___pip_5160_1_97___block_40_dt_z = _q___pip_5160_1_97___block_40_dt_z;
_d___pip_5160_1_98___block_40_dt_z = _q___pip_5160_1_98___block_40_dt_z;
_d___pip_5160_1_99___block_40_dt_z = _q___pip_5160_1_99___block_40_dt_z;
_d___pip_5160_1_100___block_40_dt_z = _q___pip_5160_1_100___block_40_dt_z;
_d___pip_5160_1_101___block_40_dt_z = _q___pip_5160_1_101___block_40_dt_z;
_d___pip_5160_1_102___block_40_dt_z = _q___pip_5160_1_102___block_40_dt_z;
_d___pip_5160_1_103___block_40_dt_z = _q___pip_5160_1_103___block_40_dt_z;
_d___pip_5160_1_104___block_40_dt_z = _q___pip_5160_1_104___block_40_dt_z;
_d___pip_5160_1_105___block_40_dt_z = _q___pip_5160_1_105___block_40_dt_z;
_d___pip_5160_1_106___block_40_dt_z = _q___pip_5160_1_106___block_40_dt_z;
_d___pip_5160_1_107___block_40_dt_z = _q___pip_5160_1_107___block_40_dt_z;
_d___pip_5160_1_108___block_40_dt_z = _q___pip_5160_1_108___block_40_dt_z;
_d___pip_5160_1_109___block_40_dt_z = _q___pip_5160_1_109___block_40_dt_z;
_d___pip_5160_1_110___block_40_dt_z = _q___pip_5160_1_110___block_40_dt_z;
_d___pip_5160_1_111___block_40_dt_z = _q___pip_5160_1_111___block_40_dt_z;
_d___pip_5160_1_112___block_40_dt_z = _q___pip_5160_1_112___block_40_dt_z;
_d___pip_5160_1_113___block_40_dt_z = _q___pip_5160_1_113___block_40_dt_z;
_d___pip_5160_1_114___block_40_dt_z = _q___pip_5160_1_114___block_40_dt_z;
_d___pip_5160_1_115___block_40_dt_z = _q___pip_5160_1_115___block_40_dt_z;
_d___pip_5160_1_116___block_40_dt_z = _q___pip_5160_1_116___block_40_dt_z;
_d___pip_5160_1_117___block_40_dt_z = _q___pip_5160_1_117___block_40_dt_z;
_d___pip_5160_1_118___block_40_dt_z = _q___pip_5160_1_118___block_40_dt_z;
_d___pip_5160_1_119___block_40_dt_z = _q___pip_5160_1_119___block_40_dt_z;
_d___pip_5160_1_120___block_40_dt_z = _q___pip_5160_1_120___block_40_dt_z;
_d___pip_5160_1_121___block_40_dt_z = _q___pip_5160_1_121___block_40_dt_z;
_d___pip_5160_1_122___block_40_dt_z = _q___pip_5160_1_122___block_40_dt_z;
_d___pip_5160_1_123___block_40_dt_z = _q___pip_5160_1_123___block_40_dt_z;
_d___pip_5160_1_124___block_40_dt_z = _q___pip_5160_1_124___block_40_dt_z;
_d___pip_5160_1_125___block_40_dt_z = _q___pip_5160_1_125___block_40_dt_z;
_d___pip_5160_1_126___block_40_dt_z = _q___pip_5160_1_126___block_40_dt_z;
_d___pip_5160_1_127___block_40_dt_z = _q___pip_5160_1_127___block_40_dt_z;
_d___pip_5160_1_128___block_40_dt_z = _q___pip_5160_1_128___block_40_dt_z;
_d___pip_5160_1_129___block_40_dt_z = _q___pip_5160_1_129___block_40_dt_z;
_d___pip_5160_1_130___block_40_dt_z = _q___pip_5160_1_130___block_40_dt_z;
_d___pip_5160_1_131___block_40_dt_z = _q___pip_5160_1_131___block_40_dt_z;
_d___pip_5160_1_132___block_40_dt_z = _q___pip_5160_1_132___block_40_dt_z;
_d___pip_5160_1_133___block_40_dt_z = _q___pip_5160_1_133___block_40_dt_z;
_d___pip_5160_1_134___block_40_dt_z = _q___pip_5160_1_134___block_40_dt_z;
_d___pip_5160_1_4___stage___block_26_brd_x = _q___pip_5160_1_4___stage___block_26_brd_x;
_d___pip_5160_1_5___stage___block_26_brd_x = _q___pip_5160_1_5___stage___block_26_brd_x;
_d___pip_5160_1_6___stage___block_26_brd_x = _q___pip_5160_1_6___stage___block_26_brd_x;
_d___pip_5160_1_4___stage___block_26_brd_y = _q___pip_5160_1_4___stage___block_26_brd_y;
_d___pip_5160_1_5___stage___block_26_brd_y = _q___pip_5160_1_5___stage___block_26_brd_y;
_d___pip_5160_1_6___stage___block_26_brd_y = _q___pip_5160_1_6___stage___block_26_brd_y;
_d___pip_5160_1_4___stage___block_26_brd_z = _q___pip_5160_1_4___stage___block_26_brd_z;
_d___pip_5160_1_5___stage___block_26_brd_z = _q___pip_5160_1_5___stage___block_26_brd_z;
_d___pip_5160_1_6___stage___block_26_brd_z = _q___pip_5160_1_6___stage___block_26_brd_z;
_d___pip_5160_1_4___stage___block_26_rd_x = _q___pip_5160_1_4___stage___block_26_rd_x;
_d___pip_5160_1_5___stage___block_26_rd_x = _q___pip_5160_1_5___stage___block_26_rd_x;
_d___pip_5160_1_4___stage___block_26_rd_y = _q___pip_5160_1_4___stage___block_26_rd_y;
_d___pip_5160_1_5___stage___block_26_rd_y = _q___pip_5160_1_5___stage___block_26_rd_y;
_d___pip_5160_1_4___stage___block_26_rd_z = _q___pip_5160_1_4___stage___block_26_rd_z;
_d___pip_5160_1_5___stage___block_26_rd_z = _q___pip_5160_1_5___stage___block_26_rd_z;
_d___pip_5160_1_4___stage___block_26_s_x = _q___pip_5160_1_4___stage___block_26_s_x;
_d___pip_5160_1_5___stage___block_26_s_x = _q___pip_5160_1_5___stage___block_26_s_x;
_d___pip_5160_1_6___stage___block_26_s_x = _q___pip_5160_1_6___stage___block_26_s_x;
_d___pip_5160_1_7___stage___block_26_s_x = _q___pip_5160_1_7___stage___block_26_s_x;
_d___pip_5160_1_8___stage___block_26_s_x = _q___pip_5160_1_8___stage___block_26_s_x;
_d___pip_5160_1_9___stage___block_26_s_x = _q___pip_5160_1_9___stage___block_26_s_x;
_d___pip_5160_1_10___stage___block_26_s_x = _q___pip_5160_1_10___stage___block_26_s_x;
_d___pip_5160_1_11___stage___block_26_s_x = _q___pip_5160_1_11___stage___block_26_s_x;
_d___pip_5160_1_12___stage___block_26_s_x = _q___pip_5160_1_12___stage___block_26_s_x;
_d___pip_5160_1_13___stage___block_26_s_x = _q___pip_5160_1_13___stage___block_26_s_x;
_d___pip_5160_1_14___stage___block_26_s_x = _q___pip_5160_1_14___stage___block_26_s_x;
_d___pip_5160_1_15___stage___block_26_s_x = _q___pip_5160_1_15___stage___block_26_s_x;
_d___pip_5160_1_16___stage___block_26_s_x = _q___pip_5160_1_16___stage___block_26_s_x;
_d___pip_5160_1_17___stage___block_26_s_x = _q___pip_5160_1_17___stage___block_26_s_x;
_d___pip_5160_1_18___stage___block_26_s_x = _q___pip_5160_1_18___stage___block_26_s_x;
_d___pip_5160_1_19___stage___block_26_s_x = _q___pip_5160_1_19___stage___block_26_s_x;
_d___pip_5160_1_20___stage___block_26_s_x = _q___pip_5160_1_20___stage___block_26_s_x;
_d___pip_5160_1_21___stage___block_26_s_x = _q___pip_5160_1_21___stage___block_26_s_x;
_d___pip_5160_1_22___stage___block_26_s_x = _q___pip_5160_1_22___stage___block_26_s_x;
_d___pip_5160_1_23___stage___block_26_s_x = _q___pip_5160_1_23___stage___block_26_s_x;
_d___pip_5160_1_24___stage___block_26_s_x = _q___pip_5160_1_24___stage___block_26_s_x;
_d___pip_5160_1_25___stage___block_26_s_x = _q___pip_5160_1_25___stage___block_26_s_x;
_d___pip_5160_1_26___stage___block_26_s_x = _q___pip_5160_1_26___stage___block_26_s_x;
_d___pip_5160_1_27___stage___block_26_s_x = _q___pip_5160_1_27___stage___block_26_s_x;
_d___pip_5160_1_28___stage___block_26_s_x = _q___pip_5160_1_28___stage___block_26_s_x;
_d___pip_5160_1_29___stage___block_26_s_x = _q___pip_5160_1_29___stage___block_26_s_x;
_d___pip_5160_1_30___stage___block_26_s_x = _q___pip_5160_1_30___stage___block_26_s_x;
_d___pip_5160_1_31___stage___block_26_s_x = _q___pip_5160_1_31___stage___block_26_s_x;
_d___pip_5160_1_32___stage___block_26_s_x = _q___pip_5160_1_32___stage___block_26_s_x;
_d___pip_5160_1_33___stage___block_26_s_x = _q___pip_5160_1_33___stage___block_26_s_x;
_d___pip_5160_1_34___stage___block_26_s_x = _q___pip_5160_1_34___stage___block_26_s_x;
_d___pip_5160_1_35___stage___block_26_s_x = _q___pip_5160_1_35___stage___block_26_s_x;
_d___pip_5160_1_36___stage___block_26_s_x = _q___pip_5160_1_36___stage___block_26_s_x;
_d___pip_5160_1_37___stage___block_26_s_x = _q___pip_5160_1_37___stage___block_26_s_x;
_d___pip_5160_1_38___stage___block_26_s_x = _q___pip_5160_1_38___stage___block_26_s_x;
_d___pip_5160_1_39___stage___block_26_s_x = _q___pip_5160_1_39___stage___block_26_s_x;
_d___pip_5160_1_40___stage___block_26_s_x = _q___pip_5160_1_40___stage___block_26_s_x;
_d___pip_5160_1_41___stage___block_26_s_x = _q___pip_5160_1_41___stage___block_26_s_x;
_d___pip_5160_1_42___stage___block_26_s_x = _q___pip_5160_1_42___stage___block_26_s_x;
_d___pip_5160_1_43___stage___block_26_s_x = _q___pip_5160_1_43___stage___block_26_s_x;
_d___pip_5160_1_44___stage___block_26_s_x = _q___pip_5160_1_44___stage___block_26_s_x;
_d___pip_5160_1_45___stage___block_26_s_x = _q___pip_5160_1_45___stage___block_26_s_x;
_d___pip_5160_1_46___stage___block_26_s_x = _q___pip_5160_1_46___stage___block_26_s_x;
_d___pip_5160_1_47___stage___block_26_s_x = _q___pip_5160_1_47___stage___block_26_s_x;
_d___pip_5160_1_48___stage___block_26_s_x = _q___pip_5160_1_48___stage___block_26_s_x;
_d___pip_5160_1_49___stage___block_26_s_x = _q___pip_5160_1_49___stage___block_26_s_x;
_d___pip_5160_1_50___stage___block_26_s_x = _q___pip_5160_1_50___stage___block_26_s_x;
_d___pip_5160_1_51___stage___block_26_s_x = _q___pip_5160_1_51___stage___block_26_s_x;
_d___pip_5160_1_52___stage___block_26_s_x = _q___pip_5160_1_52___stage___block_26_s_x;
_d___pip_5160_1_53___stage___block_26_s_x = _q___pip_5160_1_53___stage___block_26_s_x;
_d___pip_5160_1_54___stage___block_26_s_x = _q___pip_5160_1_54___stage___block_26_s_x;
_d___pip_5160_1_55___stage___block_26_s_x = _q___pip_5160_1_55___stage___block_26_s_x;
_d___pip_5160_1_56___stage___block_26_s_x = _q___pip_5160_1_56___stage___block_26_s_x;
_d___pip_5160_1_57___stage___block_26_s_x = _q___pip_5160_1_57___stage___block_26_s_x;
_d___pip_5160_1_58___stage___block_26_s_x = _q___pip_5160_1_58___stage___block_26_s_x;
_d___pip_5160_1_59___stage___block_26_s_x = _q___pip_5160_1_59___stage___block_26_s_x;
_d___pip_5160_1_60___stage___block_26_s_x = _q___pip_5160_1_60___stage___block_26_s_x;
_d___pip_5160_1_61___stage___block_26_s_x = _q___pip_5160_1_61___stage___block_26_s_x;
_d___pip_5160_1_62___stage___block_26_s_x = _q___pip_5160_1_62___stage___block_26_s_x;
_d___pip_5160_1_63___stage___block_26_s_x = _q___pip_5160_1_63___stage___block_26_s_x;
_d___pip_5160_1_64___stage___block_26_s_x = _q___pip_5160_1_64___stage___block_26_s_x;
_d___pip_5160_1_65___stage___block_26_s_x = _q___pip_5160_1_65___stage___block_26_s_x;
_d___pip_5160_1_66___stage___block_26_s_x = _q___pip_5160_1_66___stage___block_26_s_x;
_d___pip_5160_1_67___stage___block_26_s_x = _q___pip_5160_1_67___stage___block_26_s_x;
_d___pip_5160_1_68___stage___block_26_s_x = _q___pip_5160_1_68___stage___block_26_s_x;
_d___pip_5160_1_69___stage___block_26_s_x = _q___pip_5160_1_69___stage___block_26_s_x;
_d___pip_5160_1_70___stage___block_26_s_x = _q___pip_5160_1_70___stage___block_26_s_x;
_d___pip_5160_1_71___stage___block_26_s_x = _q___pip_5160_1_71___stage___block_26_s_x;
_d___pip_5160_1_72___stage___block_26_s_x = _q___pip_5160_1_72___stage___block_26_s_x;
_d___pip_5160_1_73___stage___block_26_s_x = _q___pip_5160_1_73___stage___block_26_s_x;
_d___pip_5160_1_74___stage___block_26_s_x = _q___pip_5160_1_74___stage___block_26_s_x;
_d___pip_5160_1_75___stage___block_26_s_x = _q___pip_5160_1_75___stage___block_26_s_x;
_d___pip_5160_1_76___stage___block_26_s_x = _q___pip_5160_1_76___stage___block_26_s_x;
_d___pip_5160_1_77___stage___block_26_s_x = _q___pip_5160_1_77___stage___block_26_s_x;
_d___pip_5160_1_78___stage___block_26_s_x = _q___pip_5160_1_78___stage___block_26_s_x;
_d___pip_5160_1_79___stage___block_26_s_x = _q___pip_5160_1_79___stage___block_26_s_x;
_d___pip_5160_1_80___stage___block_26_s_x = _q___pip_5160_1_80___stage___block_26_s_x;
_d___pip_5160_1_81___stage___block_26_s_x = _q___pip_5160_1_81___stage___block_26_s_x;
_d___pip_5160_1_82___stage___block_26_s_x = _q___pip_5160_1_82___stage___block_26_s_x;
_d___pip_5160_1_83___stage___block_26_s_x = _q___pip_5160_1_83___stage___block_26_s_x;
_d___pip_5160_1_84___stage___block_26_s_x = _q___pip_5160_1_84___stage___block_26_s_x;
_d___pip_5160_1_85___stage___block_26_s_x = _q___pip_5160_1_85___stage___block_26_s_x;
_d___pip_5160_1_86___stage___block_26_s_x = _q___pip_5160_1_86___stage___block_26_s_x;
_d___pip_5160_1_87___stage___block_26_s_x = _q___pip_5160_1_87___stage___block_26_s_x;
_d___pip_5160_1_88___stage___block_26_s_x = _q___pip_5160_1_88___stage___block_26_s_x;
_d___pip_5160_1_89___stage___block_26_s_x = _q___pip_5160_1_89___stage___block_26_s_x;
_d___pip_5160_1_90___stage___block_26_s_x = _q___pip_5160_1_90___stage___block_26_s_x;
_d___pip_5160_1_91___stage___block_26_s_x = _q___pip_5160_1_91___stage___block_26_s_x;
_d___pip_5160_1_92___stage___block_26_s_x = _q___pip_5160_1_92___stage___block_26_s_x;
_d___pip_5160_1_93___stage___block_26_s_x = _q___pip_5160_1_93___stage___block_26_s_x;
_d___pip_5160_1_94___stage___block_26_s_x = _q___pip_5160_1_94___stage___block_26_s_x;
_d___pip_5160_1_95___stage___block_26_s_x = _q___pip_5160_1_95___stage___block_26_s_x;
_d___pip_5160_1_96___stage___block_26_s_x = _q___pip_5160_1_96___stage___block_26_s_x;
_d___pip_5160_1_97___stage___block_26_s_x = _q___pip_5160_1_97___stage___block_26_s_x;
_d___pip_5160_1_98___stage___block_26_s_x = _q___pip_5160_1_98___stage___block_26_s_x;
_d___pip_5160_1_99___stage___block_26_s_x = _q___pip_5160_1_99___stage___block_26_s_x;
_d___pip_5160_1_100___stage___block_26_s_x = _q___pip_5160_1_100___stage___block_26_s_x;
_d___pip_5160_1_101___stage___block_26_s_x = _q___pip_5160_1_101___stage___block_26_s_x;
_d___pip_5160_1_102___stage___block_26_s_x = _q___pip_5160_1_102___stage___block_26_s_x;
_d___pip_5160_1_103___stage___block_26_s_x = _q___pip_5160_1_103___stage___block_26_s_x;
_d___pip_5160_1_104___stage___block_26_s_x = _q___pip_5160_1_104___stage___block_26_s_x;
_d___pip_5160_1_105___stage___block_26_s_x = _q___pip_5160_1_105___stage___block_26_s_x;
_d___pip_5160_1_106___stage___block_26_s_x = _q___pip_5160_1_106___stage___block_26_s_x;
_d___pip_5160_1_107___stage___block_26_s_x = _q___pip_5160_1_107___stage___block_26_s_x;
_d___pip_5160_1_108___stage___block_26_s_x = _q___pip_5160_1_108___stage___block_26_s_x;
_d___pip_5160_1_109___stage___block_26_s_x = _q___pip_5160_1_109___stage___block_26_s_x;
_d___pip_5160_1_110___stage___block_26_s_x = _q___pip_5160_1_110___stage___block_26_s_x;
_d___pip_5160_1_111___stage___block_26_s_x = _q___pip_5160_1_111___stage___block_26_s_x;
_d___pip_5160_1_112___stage___block_26_s_x = _q___pip_5160_1_112___stage___block_26_s_x;
_d___pip_5160_1_113___stage___block_26_s_x = _q___pip_5160_1_113___stage___block_26_s_x;
_d___pip_5160_1_114___stage___block_26_s_x = _q___pip_5160_1_114___stage___block_26_s_x;
_d___pip_5160_1_115___stage___block_26_s_x = _q___pip_5160_1_115___stage___block_26_s_x;
_d___pip_5160_1_116___stage___block_26_s_x = _q___pip_5160_1_116___stage___block_26_s_x;
_d___pip_5160_1_117___stage___block_26_s_x = _q___pip_5160_1_117___stage___block_26_s_x;
_d___pip_5160_1_118___stage___block_26_s_x = _q___pip_5160_1_118___stage___block_26_s_x;
_d___pip_5160_1_119___stage___block_26_s_x = _q___pip_5160_1_119___stage___block_26_s_x;
_d___pip_5160_1_120___stage___block_26_s_x = _q___pip_5160_1_120___stage___block_26_s_x;
_d___pip_5160_1_121___stage___block_26_s_x = _q___pip_5160_1_121___stage___block_26_s_x;
_d___pip_5160_1_122___stage___block_26_s_x = _q___pip_5160_1_122___stage___block_26_s_x;
_d___pip_5160_1_123___stage___block_26_s_x = _q___pip_5160_1_123___stage___block_26_s_x;
_d___pip_5160_1_124___stage___block_26_s_x = _q___pip_5160_1_124___stage___block_26_s_x;
_d___pip_5160_1_125___stage___block_26_s_x = _q___pip_5160_1_125___stage___block_26_s_x;
_d___pip_5160_1_126___stage___block_26_s_x = _q___pip_5160_1_126___stage___block_26_s_x;
_d___pip_5160_1_127___stage___block_26_s_x = _q___pip_5160_1_127___stage___block_26_s_x;
_d___pip_5160_1_128___stage___block_26_s_x = _q___pip_5160_1_128___stage___block_26_s_x;
_d___pip_5160_1_129___stage___block_26_s_x = _q___pip_5160_1_129___stage___block_26_s_x;
_d___pip_5160_1_130___stage___block_26_s_x = _q___pip_5160_1_130___stage___block_26_s_x;
_d___pip_5160_1_131___stage___block_26_s_x = _q___pip_5160_1_131___stage___block_26_s_x;
_d___pip_5160_1_132___stage___block_26_s_x = _q___pip_5160_1_132___stage___block_26_s_x;
_d___pip_5160_1_133___stage___block_26_s_x = _q___pip_5160_1_133___stage___block_26_s_x;
_d___pip_5160_1_134___stage___block_26_s_x = _q___pip_5160_1_134___stage___block_26_s_x;
_d___pip_5160_1_4___stage___block_26_s_y = _q___pip_5160_1_4___stage___block_26_s_y;
_d___pip_5160_1_5___stage___block_26_s_y = _q___pip_5160_1_5___stage___block_26_s_y;
_d___pip_5160_1_6___stage___block_26_s_y = _q___pip_5160_1_6___stage___block_26_s_y;
_d___pip_5160_1_7___stage___block_26_s_y = _q___pip_5160_1_7___stage___block_26_s_y;
_d___pip_5160_1_8___stage___block_26_s_y = _q___pip_5160_1_8___stage___block_26_s_y;
_d___pip_5160_1_9___stage___block_26_s_y = _q___pip_5160_1_9___stage___block_26_s_y;
_d___pip_5160_1_10___stage___block_26_s_y = _q___pip_5160_1_10___stage___block_26_s_y;
_d___pip_5160_1_11___stage___block_26_s_y = _q___pip_5160_1_11___stage___block_26_s_y;
_d___pip_5160_1_12___stage___block_26_s_y = _q___pip_5160_1_12___stage___block_26_s_y;
_d___pip_5160_1_13___stage___block_26_s_y = _q___pip_5160_1_13___stage___block_26_s_y;
_d___pip_5160_1_14___stage___block_26_s_y = _q___pip_5160_1_14___stage___block_26_s_y;
_d___pip_5160_1_15___stage___block_26_s_y = _q___pip_5160_1_15___stage___block_26_s_y;
_d___pip_5160_1_16___stage___block_26_s_y = _q___pip_5160_1_16___stage___block_26_s_y;
_d___pip_5160_1_17___stage___block_26_s_y = _q___pip_5160_1_17___stage___block_26_s_y;
_d___pip_5160_1_18___stage___block_26_s_y = _q___pip_5160_1_18___stage___block_26_s_y;
_d___pip_5160_1_19___stage___block_26_s_y = _q___pip_5160_1_19___stage___block_26_s_y;
_d___pip_5160_1_20___stage___block_26_s_y = _q___pip_5160_1_20___stage___block_26_s_y;
_d___pip_5160_1_21___stage___block_26_s_y = _q___pip_5160_1_21___stage___block_26_s_y;
_d___pip_5160_1_22___stage___block_26_s_y = _q___pip_5160_1_22___stage___block_26_s_y;
_d___pip_5160_1_23___stage___block_26_s_y = _q___pip_5160_1_23___stage___block_26_s_y;
_d___pip_5160_1_24___stage___block_26_s_y = _q___pip_5160_1_24___stage___block_26_s_y;
_d___pip_5160_1_25___stage___block_26_s_y = _q___pip_5160_1_25___stage___block_26_s_y;
_d___pip_5160_1_26___stage___block_26_s_y = _q___pip_5160_1_26___stage___block_26_s_y;
_d___pip_5160_1_27___stage___block_26_s_y = _q___pip_5160_1_27___stage___block_26_s_y;
_d___pip_5160_1_28___stage___block_26_s_y = _q___pip_5160_1_28___stage___block_26_s_y;
_d___pip_5160_1_29___stage___block_26_s_y = _q___pip_5160_1_29___stage___block_26_s_y;
_d___pip_5160_1_30___stage___block_26_s_y = _q___pip_5160_1_30___stage___block_26_s_y;
_d___pip_5160_1_31___stage___block_26_s_y = _q___pip_5160_1_31___stage___block_26_s_y;
_d___pip_5160_1_32___stage___block_26_s_y = _q___pip_5160_1_32___stage___block_26_s_y;
_d___pip_5160_1_33___stage___block_26_s_y = _q___pip_5160_1_33___stage___block_26_s_y;
_d___pip_5160_1_34___stage___block_26_s_y = _q___pip_5160_1_34___stage___block_26_s_y;
_d___pip_5160_1_35___stage___block_26_s_y = _q___pip_5160_1_35___stage___block_26_s_y;
_d___pip_5160_1_36___stage___block_26_s_y = _q___pip_5160_1_36___stage___block_26_s_y;
_d___pip_5160_1_37___stage___block_26_s_y = _q___pip_5160_1_37___stage___block_26_s_y;
_d___pip_5160_1_38___stage___block_26_s_y = _q___pip_5160_1_38___stage___block_26_s_y;
_d___pip_5160_1_39___stage___block_26_s_y = _q___pip_5160_1_39___stage___block_26_s_y;
_d___pip_5160_1_40___stage___block_26_s_y = _q___pip_5160_1_40___stage___block_26_s_y;
_d___pip_5160_1_41___stage___block_26_s_y = _q___pip_5160_1_41___stage___block_26_s_y;
_d___pip_5160_1_42___stage___block_26_s_y = _q___pip_5160_1_42___stage___block_26_s_y;
_d___pip_5160_1_43___stage___block_26_s_y = _q___pip_5160_1_43___stage___block_26_s_y;
_d___pip_5160_1_44___stage___block_26_s_y = _q___pip_5160_1_44___stage___block_26_s_y;
_d___pip_5160_1_45___stage___block_26_s_y = _q___pip_5160_1_45___stage___block_26_s_y;
_d___pip_5160_1_46___stage___block_26_s_y = _q___pip_5160_1_46___stage___block_26_s_y;
_d___pip_5160_1_47___stage___block_26_s_y = _q___pip_5160_1_47___stage___block_26_s_y;
_d___pip_5160_1_48___stage___block_26_s_y = _q___pip_5160_1_48___stage___block_26_s_y;
_d___pip_5160_1_49___stage___block_26_s_y = _q___pip_5160_1_49___stage___block_26_s_y;
_d___pip_5160_1_50___stage___block_26_s_y = _q___pip_5160_1_50___stage___block_26_s_y;
_d___pip_5160_1_51___stage___block_26_s_y = _q___pip_5160_1_51___stage___block_26_s_y;
_d___pip_5160_1_52___stage___block_26_s_y = _q___pip_5160_1_52___stage___block_26_s_y;
_d___pip_5160_1_53___stage___block_26_s_y = _q___pip_5160_1_53___stage___block_26_s_y;
_d___pip_5160_1_54___stage___block_26_s_y = _q___pip_5160_1_54___stage___block_26_s_y;
_d___pip_5160_1_55___stage___block_26_s_y = _q___pip_5160_1_55___stage___block_26_s_y;
_d___pip_5160_1_56___stage___block_26_s_y = _q___pip_5160_1_56___stage___block_26_s_y;
_d___pip_5160_1_57___stage___block_26_s_y = _q___pip_5160_1_57___stage___block_26_s_y;
_d___pip_5160_1_58___stage___block_26_s_y = _q___pip_5160_1_58___stage___block_26_s_y;
_d___pip_5160_1_59___stage___block_26_s_y = _q___pip_5160_1_59___stage___block_26_s_y;
_d___pip_5160_1_60___stage___block_26_s_y = _q___pip_5160_1_60___stage___block_26_s_y;
_d___pip_5160_1_61___stage___block_26_s_y = _q___pip_5160_1_61___stage___block_26_s_y;
_d___pip_5160_1_62___stage___block_26_s_y = _q___pip_5160_1_62___stage___block_26_s_y;
_d___pip_5160_1_63___stage___block_26_s_y = _q___pip_5160_1_63___stage___block_26_s_y;
_d___pip_5160_1_64___stage___block_26_s_y = _q___pip_5160_1_64___stage___block_26_s_y;
_d___pip_5160_1_65___stage___block_26_s_y = _q___pip_5160_1_65___stage___block_26_s_y;
_d___pip_5160_1_66___stage___block_26_s_y = _q___pip_5160_1_66___stage___block_26_s_y;
_d___pip_5160_1_67___stage___block_26_s_y = _q___pip_5160_1_67___stage___block_26_s_y;
_d___pip_5160_1_68___stage___block_26_s_y = _q___pip_5160_1_68___stage___block_26_s_y;
_d___pip_5160_1_69___stage___block_26_s_y = _q___pip_5160_1_69___stage___block_26_s_y;
_d___pip_5160_1_70___stage___block_26_s_y = _q___pip_5160_1_70___stage___block_26_s_y;
_d___pip_5160_1_71___stage___block_26_s_y = _q___pip_5160_1_71___stage___block_26_s_y;
_d___pip_5160_1_72___stage___block_26_s_y = _q___pip_5160_1_72___stage___block_26_s_y;
_d___pip_5160_1_73___stage___block_26_s_y = _q___pip_5160_1_73___stage___block_26_s_y;
_d___pip_5160_1_74___stage___block_26_s_y = _q___pip_5160_1_74___stage___block_26_s_y;
_d___pip_5160_1_75___stage___block_26_s_y = _q___pip_5160_1_75___stage___block_26_s_y;
_d___pip_5160_1_76___stage___block_26_s_y = _q___pip_5160_1_76___stage___block_26_s_y;
_d___pip_5160_1_77___stage___block_26_s_y = _q___pip_5160_1_77___stage___block_26_s_y;
_d___pip_5160_1_78___stage___block_26_s_y = _q___pip_5160_1_78___stage___block_26_s_y;
_d___pip_5160_1_79___stage___block_26_s_y = _q___pip_5160_1_79___stage___block_26_s_y;
_d___pip_5160_1_80___stage___block_26_s_y = _q___pip_5160_1_80___stage___block_26_s_y;
_d___pip_5160_1_81___stage___block_26_s_y = _q___pip_5160_1_81___stage___block_26_s_y;
_d___pip_5160_1_82___stage___block_26_s_y = _q___pip_5160_1_82___stage___block_26_s_y;
_d___pip_5160_1_83___stage___block_26_s_y = _q___pip_5160_1_83___stage___block_26_s_y;
_d___pip_5160_1_84___stage___block_26_s_y = _q___pip_5160_1_84___stage___block_26_s_y;
_d___pip_5160_1_85___stage___block_26_s_y = _q___pip_5160_1_85___stage___block_26_s_y;
_d___pip_5160_1_86___stage___block_26_s_y = _q___pip_5160_1_86___stage___block_26_s_y;
_d___pip_5160_1_87___stage___block_26_s_y = _q___pip_5160_1_87___stage___block_26_s_y;
_d___pip_5160_1_88___stage___block_26_s_y = _q___pip_5160_1_88___stage___block_26_s_y;
_d___pip_5160_1_89___stage___block_26_s_y = _q___pip_5160_1_89___stage___block_26_s_y;
_d___pip_5160_1_90___stage___block_26_s_y = _q___pip_5160_1_90___stage___block_26_s_y;
_d___pip_5160_1_91___stage___block_26_s_y = _q___pip_5160_1_91___stage___block_26_s_y;
_d___pip_5160_1_92___stage___block_26_s_y = _q___pip_5160_1_92___stage___block_26_s_y;
_d___pip_5160_1_93___stage___block_26_s_y = _q___pip_5160_1_93___stage___block_26_s_y;
_d___pip_5160_1_94___stage___block_26_s_y = _q___pip_5160_1_94___stage___block_26_s_y;
_d___pip_5160_1_95___stage___block_26_s_y = _q___pip_5160_1_95___stage___block_26_s_y;
_d___pip_5160_1_96___stage___block_26_s_y = _q___pip_5160_1_96___stage___block_26_s_y;
_d___pip_5160_1_97___stage___block_26_s_y = _q___pip_5160_1_97___stage___block_26_s_y;
_d___pip_5160_1_98___stage___block_26_s_y = _q___pip_5160_1_98___stage___block_26_s_y;
_d___pip_5160_1_99___stage___block_26_s_y = _q___pip_5160_1_99___stage___block_26_s_y;
_d___pip_5160_1_100___stage___block_26_s_y = _q___pip_5160_1_100___stage___block_26_s_y;
_d___pip_5160_1_101___stage___block_26_s_y = _q___pip_5160_1_101___stage___block_26_s_y;
_d___pip_5160_1_102___stage___block_26_s_y = _q___pip_5160_1_102___stage___block_26_s_y;
_d___pip_5160_1_103___stage___block_26_s_y = _q___pip_5160_1_103___stage___block_26_s_y;
_d___pip_5160_1_104___stage___block_26_s_y = _q___pip_5160_1_104___stage___block_26_s_y;
_d___pip_5160_1_105___stage___block_26_s_y = _q___pip_5160_1_105___stage___block_26_s_y;
_d___pip_5160_1_106___stage___block_26_s_y = _q___pip_5160_1_106___stage___block_26_s_y;
_d___pip_5160_1_107___stage___block_26_s_y = _q___pip_5160_1_107___stage___block_26_s_y;
_d___pip_5160_1_108___stage___block_26_s_y = _q___pip_5160_1_108___stage___block_26_s_y;
_d___pip_5160_1_109___stage___block_26_s_y = _q___pip_5160_1_109___stage___block_26_s_y;
_d___pip_5160_1_110___stage___block_26_s_y = _q___pip_5160_1_110___stage___block_26_s_y;
_d___pip_5160_1_111___stage___block_26_s_y = _q___pip_5160_1_111___stage___block_26_s_y;
_d___pip_5160_1_112___stage___block_26_s_y = _q___pip_5160_1_112___stage___block_26_s_y;
_d___pip_5160_1_113___stage___block_26_s_y = _q___pip_5160_1_113___stage___block_26_s_y;
_d___pip_5160_1_114___stage___block_26_s_y = _q___pip_5160_1_114___stage___block_26_s_y;
_d___pip_5160_1_115___stage___block_26_s_y = _q___pip_5160_1_115___stage___block_26_s_y;
_d___pip_5160_1_116___stage___block_26_s_y = _q___pip_5160_1_116___stage___block_26_s_y;
_d___pip_5160_1_117___stage___block_26_s_y = _q___pip_5160_1_117___stage___block_26_s_y;
_d___pip_5160_1_118___stage___block_26_s_y = _q___pip_5160_1_118___stage___block_26_s_y;
_d___pip_5160_1_119___stage___block_26_s_y = _q___pip_5160_1_119___stage___block_26_s_y;
_d___pip_5160_1_120___stage___block_26_s_y = _q___pip_5160_1_120___stage___block_26_s_y;
_d___pip_5160_1_121___stage___block_26_s_y = _q___pip_5160_1_121___stage___block_26_s_y;
_d___pip_5160_1_122___stage___block_26_s_y = _q___pip_5160_1_122___stage___block_26_s_y;
_d___pip_5160_1_123___stage___block_26_s_y = _q___pip_5160_1_123___stage___block_26_s_y;
_d___pip_5160_1_124___stage___block_26_s_y = _q___pip_5160_1_124___stage___block_26_s_y;
_d___pip_5160_1_125___stage___block_26_s_y = _q___pip_5160_1_125___stage___block_26_s_y;
_d___pip_5160_1_126___stage___block_26_s_y = _q___pip_5160_1_126___stage___block_26_s_y;
_d___pip_5160_1_127___stage___block_26_s_y = _q___pip_5160_1_127___stage___block_26_s_y;
_d___pip_5160_1_128___stage___block_26_s_y = _q___pip_5160_1_128___stage___block_26_s_y;
_d___pip_5160_1_129___stage___block_26_s_y = _q___pip_5160_1_129___stage___block_26_s_y;
_d___pip_5160_1_130___stage___block_26_s_y = _q___pip_5160_1_130___stage___block_26_s_y;
_d___pip_5160_1_131___stage___block_26_s_y = _q___pip_5160_1_131___stage___block_26_s_y;
_d___pip_5160_1_132___stage___block_26_s_y = _q___pip_5160_1_132___stage___block_26_s_y;
_d___pip_5160_1_133___stage___block_26_s_y = _q___pip_5160_1_133___stage___block_26_s_y;
_d___pip_5160_1_134___stage___block_26_s_y = _q___pip_5160_1_134___stage___block_26_s_y;
_d___pip_5160_1_4___stage___block_26_s_z = _q___pip_5160_1_4___stage___block_26_s_z;
_d___pip_5160_1_5___stage___block_26_s_z = _q___pip_5160_1_5___stage___block_26_s_z;
_d___pip_5160_1_6___stage___block_26_s_z = _q___pip_5160_1_6___stage___block_26_s_z;
_d___pip_5160_1_7___stage___block_26_s_z = _q___pip_5160_1_7___stage___block_26_s_z;
_d___pip_5160_1_8___stage___block_26_s_z = _q___pip_5160_1_8___stage___block_26_s_z;
_d___pip_5160_1_9___stage___block_26_s_z = _q___pip_5160_1_9___stage___block_26_s_z;
_d___pip_5160_1_10___stage___block_26_s_z = _q___pip_5160_1_10___stage___block_26_s_z;
_d___pip_5160_1_11___stage___block_26_s_z = _q___pip_5160_1_11___stage___block_26_s_z;
_d___pip_5160_1_12___stage___block_26_s_z = _q___pip_5160_1_12___stage___block_26_s_z;
_d___pip_5160_1_13___stage___block_26_s_z = _q___pip_5160_1_13___stage___block_26_s_z;
_d___pip_5160_1_14___stage___block_26_s_z = _q___pip_5160_1_14___stage___block_26_s_z;
_d___pip_5160_1_15___stage___block_26_s_z = _q___pip_5160_1_15___stage___block_26_s_z;
_d___pip_5160_1_16___stage___block_26_s_z = _q___pip_5160_1_16___stage___block_26_s_z;
_d___pip_5160_1_17___stage___block_26_s_z = _q___pip_5160_1_17___stage___block_26_s_z;
_d___pip_5160_1_18___stage___block_26_s_z = _q___pip_5160_1_18___stage___block_26_s_z;
_d___pip_5160_1_19___stage___block_26_s_z = _q___pip_5160_1_19___stage___block_26_s_z;
_d___pip_5160_1_20___stage___block_26_s_z = _q___pip_5160_1_20___stage___block_26_s_z;
_d___pip_5160_1_21___stage___block_26_s_z = _q___pip_5160_1_21___stage___block_26_s_z;
_d___pip_5160_1_22___stage___block_26_s_z = _q___pip_5160_1_22___stage___block_26_s_z;
_d___pip_5160_1_23___stage___block_26_s_z = _q___pip_5160_1_23___stage___block_26_s_z;
_d___pip_5160_1_24___stage___block_26_s_z = _q___pip_5160_1_24___stage___block_26_s_z;
_d___pip_5160_1_25___stage___block_26_s_z = _q___pip_5160_1_25___stage___block_26_s_z;
_d___pip_5160_1_26___stage___block_26_s_z = _q___pip_5160_1_26___stage___block_26_s_z;
_d___pip_5160_1_27___stage___block_26_s_z = _q___pip_5160_1_27___stage___block_26_s_z;
_d___pip_5160_1_28___stage___block_26_s_z = _q___pip_5160_1_28___stage___block_26_s_z;
_d___pip_5160_1_29___stage___block_26_s_z = _q___pip_5160_1_29___stage___block_26_s_z;
_d___pip_5160_1_30___stage___block_26_s_z = _q___pip_5160_1_30___stage___block_26_s_z;
_d___pip_5160_1_31___stage___block_26_s_z = _q___pip_5160_1_31___stage___block_26_s_z;
_d___pip_5160_1_32___stage___block_26_s_z = _q___pip_5160_1_32___stage___block_26_s_z;
_d___pip_5160_1_33___stage___block_26_s_z = _q___pip_5160_1_33___stage___block_26_s_z;
_d___pip_5160_1_34___stage___block_26_s_z = _q___pip_5160_1_34___stage___block_26_s_z;
_d___pip_5160_1_35___stage___block_26_s_z = _q___pip_5160_1_35___stage___block_26_s_z;
_d___pip_5160_1_36___stage___block_26_s_z = _q___pip_5160_1_36___stage___block_26_s_z;
_d___pip_5160_1_37___stage___block_26_s_z = _q___pip_5160_1_37___stage___block_26_s_z;
_d___pip_5160_1_38___stage___block_26_s_z = _q___pip_5160_1_38___stage___block_26_s_z;
_d___pip_5160_1_39___stage___block_26_s_z = _q___pip_5160_1_39___stage___block_26_s_z;
_d___pip_5160_1_40___stage___block_26_s_z = _q___pip_5160_1_40___stage___block_26_s_z;
_d___pip_5160_1_41___stage___block_26_s_z = _q___pip_5160_1_41___stage___block_26_s_z;
_d___pip_5160_1_42___stage___block_26_s_z = _q___pip_5160_1_42___stage___block_26_s_z;
_d___pip_5160_1_43___stage___block_26_s_z = _q___pip_5160_1_43___stage___block_26_s_z;
_d___pip_5160_1_44___stage___block_26_s_z = _q___pip_5160_1_44___stage___block_26_s_z;
_d___pip_5160_1_45___stage___block_26_s_z = _q___pip_5160_1_45___stage___block_26_s_z;
_d___pip_5160_1_46___stage___block_26_s_z = _q___pip_5160_1_46___stage___block_26_s_z;
_d___pip_5160_1_47___stage___block_26_s_z = _q___pip_5160_1_47___stage___block_26_s_z;
_d___pip_5160_1_48___stage___block_26_s_z = _q___pip_5160_1_48___stage___block_26_s_z;
_d___pip_5160_1_49___stage___block_26_s_z = _q___pip_5160_1_49___stage___block_26_s_z;
_d___pip_5160_1_50___stage___block_26_s_z = _q___pip_5160_1_50___stage___block_26_s_z;
_d___pip_5160_1_51___stage___block_26_s_z = _q___pip_5160_1_51___stage___block_26_s_z;
_d___pip_5160_1_52___stage___block_26_s_z = _q___pip_5160_1_52___stage___block_26_s_z;
_d___pip_5160_1_53___stage___block_26_s_z = _q___pip_5160_1_53___stage___block_26_s_z;
_d___pip_5160_1_54___stage___block_26_s_z = _q___pip_5160_1_54___stage___block_26_s_z;
_d___pip_5160_1_55___stage___block_26_s_z = _q___pip_5160_1_55___stage___block_26_s_z;
_d___pip_5160_1_56___stage___block_26_s_z = _q___pip_5160_1_56___stage___block_26_s_z;
_d___pip_5160_1_57___stage___block_26_s_z = _q___pip_5160_1_57___stage___block_26_s_z;
_d___pip_5160_1_58___stage___block_26_s_z = _q___pip_5160_1_58___stage___block_26_s_z;
_d___pip_5160_1_59___stage___block_26_s_z = _q___pip_5160_1_59___stage___block_26_s_z;
_d___pip_5160_1_60___stage___block_26_s_z = _q___pip_5160_1_60___stage___block_26_s_z;
_d___pip_5160_1_61___stage___block_26_s_z = _q___pip_5160_1_61___stage___block_26_s_z;
_d___pip_5160_1_62___stage___block_26_s_z = _q___pip_5160_1_62___stage___block_26_s_z;
_d___pip_5160_1_63___stage___block_26_s_z = _q___pip_5160_1_63___stage___block_26_s_z;
_d___pip_5160_1_64___stage___block_26_s_z = _q___pip_5160_1_64___stage___block_26_s_z;
_d___pip_5160_1_65___stage___block_26_s_z = _q___pip_5160_1_65___stage___block_26_s_z;
_d___pip_5160_1_66___stage___block_26_s_z = _q___pip_5160_1_66___stage___block_26_s_z;
_d___pip_5160_1_67___stage___block_26_s_z = _q___pip_5160_1_67___stage___block_26_s_z;
_d___pip_5160_1_68___stage___block_26_s_z = _q___pip_5160_1_68___stage___block_26_s_z;
_d___pip_5160_1_69___stage___block_26_s_z = _q___pip_5160_1_69___stage___block_26_s_z;
_d___pip_5160_1_70___stage___block_26_s_z = _q___pip_5160_1_70___stage___block_26_s_z;
_d___pip_5160_1_71___stage___block_26_s_z = _q___pip_5160_1_71___stage___block_26_s_z;
_d___pip_5160_1_72___stage___block_26_s_z = _q___pip_5160_1_72___stage___block_26_s_z;
_d___pip_5160_1_73___stage___block_26_s_z = _q___pip_5160_1_73___stage___block_26_s_z;
_d___pip_5160_1_74___stage___block_26_s_z = _q___pip_5160_1_74___stage___block_26_s_z;
_d___pip_5160_1_75___stage___block_26_s_z = _q___pip_5160_1_75___stage___block_26_s_z;
_d___pip_5160_1_76___stage___block_26_s_z = _q___pip_5160_1_76___stage___block_26_s_z;
_d___pip_5160_1_77___stage___block_26_s_z = _q___pip_5160_1_77___stage___block_26_s_z;
_d___pip_5160_1_78___stage___block_26_s_z = _q___pip_5160_1_78___stage___block_26_s_z;
_d___pip_5160_1_79___stage___block_26_s_z = _q___pip_5160_1_79___stage___block_26_s_z;
_d___pip_5160_1_80___stage___block_26_s_z = _q___pip_5160_1_80___stage___block_26_s_z;
_d___pip_5160_1_81___stage___block_26_s_z = _q___pip_5160_1_81___stage___block_26_s_z;
_d___pip_5160_1_82___stage___block_26_s_z = _q___pip_5160_1_82___stage___block_26_s_z;
_d___pip_5160_1_83___stage___block_26_s_z = _q___pip_5160_1_83___stage___block_26_s_z;
_d___pip_5160_1_84___stage___block_26_s_z = _q___pip_5160_1_84___stage___block_26_s_z;
_d___pip_5160_1_85___stage___block_26_s_z = _q___pip_5160_1_85___stage___block_26_s_z;
_d___pip_5160_1_86___stage___block_26_s_z = _q___pip_5160_1_86___stage___block_26_s_z;
_d___pip_5160_1_87___stage___block_26_s_z = _q___pip_5160_1_87___stage___block_26_s_z;
_d___pip_5160_1_88___stage___block_26_s_z = _q___pip_5160_1_88___stage___block_26_s_z;
_d___pip_5160_1_89___stage___block_26_s_z = _q___pip_5160_1_89___stage___block_26_s_z;
_d___pip_5160_1_90___stage___block_26_s_z = _q___pip_5160_1_90___stage___block_26_s_z;
_d___pip_5160_1_91___stage___block_26_s_z = _q___pip_5160_1_91___stage___block_26_s_z;
_d___pip_5160_1_92___stage___block_26_s_z = _q___pip_5160_1_92___stage___block_26_s_z;
_d___pip_5160_1_93___stage___block_26_s_z = _q___pip_5160_1_93___stage___block_26_s_z;
_d___pip_5160_1_94___stage___block_26_s_z = _q___pip_5160_1_94___stage___block_26_s_z;
_d___pip_5160_1_95___stage___block_26_s_z = _q___pip_5160_1_95___stage___block_26_s_z;
_d___pip_5160_1_96___stage___block_26_s_z = _q___pip_5160_1_96___stage___block_26_s_z;
_d___pip_5160_1_97___stage___block_26_s_z = _q___pip_5160_1_97___stage___block_26_s_z;
_d___pip_5160_1_98___stage___block_26_s_z = _q___pip_5160_1_98___stage___block_26_s_z;
_d___pip_5160_1_99___stage___block_26_s_z = _q___pip_5160_1_99___stage___block_26_s_z;
_d___pip_5160_1_100___stage___block_26_s_z = _q___pip_5160_1_100___stage___block_26_s_z;
_d___pip_5160_1_101___stage___block_26_s_z = _q___pip_5160_1_101___stage___block_26_s_z;
_d___pip_5160_1_102___stage___block_26_s_z = _q___pip_5160_1_102___stage___block_26_s_z;
_d___pip_5160_1_103___stage___block_26_s_z = _q___pip_5160_1_103___stage___block_26_s_z;
_d___pip_5160_1_104___stage___block_26_s_z = _q___pip_5160_1_104___stage___block_26_s_z;
_d___pip_5160_1_105___stage___block_26_s_z = _q___pip_5160_1_105___stage___block_26_s_z;
_d___pip_5160_1_106___stage___block_26_s_z = _q___pip_5160_1_106___stage___block_26_s_z;
_d___pip_5160_1_107___stage___block_26_s_z = _q___pip_5160_1_107___stage___block_26_s_z;
_d___pip_5160_1_108___stage___block_26_s_z = _q___pip_5160_1_108___stage___block_26_s_z;
_d___pip_5160_1_109___stage___block_26_s_z = _q___pip_5160_1_109___stage___block_26_s_z;
_d___pip_5160_1_110___stage___block_26_s_z = _q___pip_5160_1_110___stage___block_26_s_z;
_d___pip_5160_1_111___stage___block_26_s_z = _q___pip_5160_1_111___stage___block_26_s_z;
_d___pip_5160_1_112___stage___block_26_s_z = _q___pip_5160_1_112___stage___block_26_s_z;
_d___pip_5160_1_113___stage___block_26_s_z = _q___pip_5160_1_113___stage___block_26_s_z;
_d___pip_5160_1_114___stage___block_26_s_z = _q___pip_5160_1_114___stage___block_26_s_z;
_d___pip_5160_1_115___stage___block_26_s_z = _q___pip_5160_1_115___stage___block_26_s_z;
_d___pip_5160_1_116___stage___block_26_s_z = _q___pip_5160_1_116___stage___block_26_s_z;
_d___pip_5160_1_117___stage___block_26_s_z = _q___pip_5160_1_117___stage___block_26_s_z;
_d___pip_5160_1_118___stage___block_26_s_z = _q___pip_5160_1_118___stage___block_26_s_z;
_d___pip_5160_1_119___stage___block_26_s_z = _q___pip_5160_1_119___stage___block_26_s_z;
_d___pip_5160_1_120___stage___block_26_s_z = _q___pip_5160_1_120___stage___block_26_s_z;
_d___pip_5160_1_121___stage___block_26_s_z = _q___pip_5160_1_121___stage___block_26_s_z;
_d___pip_5160_1_122___stage___block_26_s_z = _q___pip_5160_1_122___stage___block_26_s_z;
_d___pip_5160_1_123___stage___block_26_s_z = _q___pip_5160_1_123___stage___block_26_s_z;
_d___pip_5160_1_124___stage___block_26_s_z = _q___pip_5160_1_124___stage___block_26_s_z;
_d___pip_5160_1_125___stage___block_26_s_z = _q___pip_5160_1_125___stage___block_26_s_z;
_d___pip_5160_1_126___stage___block_26_s_z = _q___pip_5160_1_126___stage___block_26_s_z;
_d___pip_5160_1_127___stage___block_26_s_z = _q___pip_5160_1_127___stage___block_26_s_z;
_d___pip_5160_1_128___stage___block_26_s_z = _q___pip_5160_1_128___stage___block_26_s_z;
_d___pip_5160_1_129___stage___block_26_s_z = _q___pip_5160_1_129___stage___block_26_s_z;
_d___pip_5160_1_130___stage___block_26_s_z = _q___pip_5160_1_130___stage___block_26_s_z;
_d___pip_5160_1_131___stage___block_26_s_z = _q___pip_5160_1_131___stage___block_26_s_z;
_d___pip_5160_1_132___stage___block_26_s_z = _q___pip_5160_1_132___stage___block_26_s_z;
_d___pip_5160_1_133___stage___block_26_s_z = _q___pip_5160_1_133___stage___block_26_s_z;
_d___pip_5160_1_134___stage___block_26_s_z = _q___pip_5160_1_134___stage___block_26_s_z;
_d___pip_5160_1_4___stage___block_26_v_x = _q___pip_5160_1_4___stage___block_26_v_x;
_d___pip_5160_1_5___stage___block_26_v_x = _q___pip_5160_1_5___stage___block_26_v_x;
_d___pip_5160_1_6___stage___block_26_v_x = _q___pip_5160_1_6___stage___block_26_v_x;
_d___pip_5160_1_7___stage___block_26_v_x = _q___pip_5160_1_7___stage___block_26_v_x;
_d___pip_5160_1_8___stage___block_26_v_x = _q___pip_5160_1_8___stage___block_26_v_x;
_d___pip_5160_1_9___stage___block_26_v_x = _q___pip_5160_1_9___stage___block_26_v_x;
_d___pip_5160_1_10___stage___block_26_v_x = _q___pip_5160_1_10___stage___block_26_v_x;
_d___pip_5160_1_11___stage___block_26_v_x = _q___pip_5160_1_11___stage___block_26_v_x;
_d___pip_5160_1_12___stage___block_26_v_x = _q___pip_5160_1_12___stage___block_26_v_x;
_d___pip_5160_1_13___stage___block_26_v_x = _q___pip_5160_1_13___stage___block_26_v_x;
_d___pip_5160_1_14___stage___block_26_v_x = _q___pip_5160_1_14___stage___block_26_v_x;
_d___pip_5160_1_15___stage___block_26_v_x = _q___pip_5160_1_15___stage___block_26_v_x;
_d___pip_5160_1_16___stage___block_26_v_x = _q___pip_5160_1_16___stage___block_26_v_x;
_d___pip_5160_1_17___stage___block_26_v_x = _q___pip_5160_1_17___stage___block_26_v_x;
_d___pip_5160_1_18___stage___block_26_v_x = _q___pip_5160_1_18___stage___block_26_v_x;
_d___pip_5160_1_19___stage___block_26_v_x = _q___pip_5160_1_19___stage___block_26_v_x;
_d___pip_5160_1_20___stage___block_26_v_x = _q___pip_5160_1_20___stage___block_26_v_x;
_d___pip_5160_1_21___stage___block_26_v_x = _q___pip_5160_1_21___stage___block_26_v_x;
_d___pip_5160_1_22___stage___block_26_v_x = _q___pip_5160_1_22___stage___block_26_v_x;
_d___pip_5160_1_23___stage___block_26_v_x = _q___pip_5160_1_23___stage___block_26_v_x;
_d___pip_5160_1_24___stage___block_26_v_x = _q___pip_5160_1_24___stage___block_26_v_x;
_d___pip_5160_1_25___stage___block_26_v_x = _q___pip_5160_1_25___stage___block_26_v_x;
_d___pip_5160_1_26___stage___block_26_v_x = _q___pip_5160_1_26___stage___block_26_v_x;
_d___pip_5160_1_27___stage___block_26_v_x = _q___pip_5160_1_27___stage___block_26_v_x;
_d___pip_5160_1_28___stage___block_26_v_x = _q___pip_5160_1_28___stage___block_26_v_x;
_d___pip_5160_1_29___stage___block_26_v_x = _q___pip_5160_1_29___stage___block_26_v_x;
_d___pip_5160_1_30___stage___block_26_v_x = _q___pip_5160_1_30___stage___block_26_v_x;
_d___pip_5160_1_31___stage___block_26_v_x = _q___pip_5160_1_31___stage___block_26_v_x;
_d___pip_5160_1_32___stage___block_26_v_x = _q___pip_5160_1_32___stage___block_26_v_x;
_d___pip_5160_1_33___stage___block_26_v_x = _q___pip_5160_1_33___stage___block_26_v_x;
_d___pip_5160_1_34___stage___block_26_v_x = _q___pip_5160_1_34___stage___block_26_v_x;
_d___pip_5160_1_35___stage___block_26_v_x = _q___pip_5160_1_35___stage___block_26_v_x;
_d___pip_5160_1_36___stage___block_26_v_x = _q___pip_5160_1_36___stage___block_26_v_x;
_d___pip_5160_1_37___stage___block_26_v_x = _q___pip_5160_1_37___stage___block_26_v_x;
_d___pip_5160_1_38___stage___block_26_v_x = _q___pip_5160_1_38___stage___block_26_v_x;
_d___pip_5160_1_39___stage___block_26_v_x = _q___pip_5160_1_39___stage___block_26_v_x;
_d___pip_5160_1_40___stage___block_26_v_x = _q___pip_5160_1_40___stage___block_26_v_x;
_d___pip_5160_1_41___stage___block_26_v_x = _q___pip_5160_1_41___stage___block_26_v_x;
_d___pip_5160_1_42___stage___block_26_v_x = _q___pip_5160_1_42___stage___block_26_v_x;
_d___pip_5160_1_43___stage___block_26_v_x = _q___pip_5160_1_43___stage___block_26_v_x;
_d___pip_5160_1_44___stage___block_26_v_x = _q___pip_5160_1_44___stage___block_26_v_x;
_d___pip_5160_1_45___stage___block_26_v_x = _q___pip_5160_1_45___stage___block_26_v_x;
_d___pip_5160_1_46___stage___block_26_v_x = _q___pip_5160_1_46___stage___block_26_v_x;
_d___pip_5160_1_47___stage___block_26_v_x = _q___pip_5160_1_47___stage___block_26_v_x;
_d___pip_5160_1_48___stage___block_26_v_x = _q___pip_5160_1_48___stage___block_26_v_x;
_d___pip_5160_1_49___stage___block_26_v_x = _q___pip_5160_1_49___stage___block_26_v_x;
_d___pip_5160_1_50___stage___block_26_v_x = _q___pip_5160_1_50___stage___block_26_v_x;
_d___pip_5160_1_51___stage___block_26_v_x = _q___pip_5160_1_51___stage___block_26_v_x;
_d___pip_5160_1_52___stage___block_26_v_x = _q___pip_5160_1_52___stage___block_26_v_x;
_d___pip_5160_1_53___stage___block_26_v_x = _q___pip_5160_1_53___stage___block_26_v_x;
_d___pip_5160_1_54___stage___block_26_v_x = _q___pip_5160_1_54___stage___block_26_v_x;
_d___pip_5160_1_55___stage___block_26_v_x = _q___pip_5160_1_55___stage___block_26_v_x;
_d___pip_5160_1_56___stage___block_26_v_x = _q___pip_5160_1_56___stage___block_26_v_x;
_d___pip_5160_1_57___stage___block_26_v_x = _q___pip_5160_1_57___stage___block_26_v_x;
_d___pip_5160_1_58___stage___block_26_v_x = _q___pip_5160_1_58___stage___block_26_v_x;
_d___pip_5160_1_59___stage___block_26_v_x = _q___pip_5160_1_59___stage___block_26_v_x;
_d___pip_5160_1_60___stage___block_26_v_x = _q___pip_5160_1_60___stage___block_26_v_x;
_d___pip_5160_1_61___stage___block_26_v_x = _q___pip_5160_1_61___stage___block_26_v_x;
_d___pip_5160_1_62___stage___block_26_v_x = _q___pip_5160_1_62___stage___block_26_v_x;
_d___pip_5160_1_63___stage___block_26_v_x = _q___pip_5160_1_63___stage___block_26_v_x;
_d___pip_5160_1_64___stage___block_26_v_x = _q___pip_5160_1_64___stage___block_26_v_x;
_d___pip_5160_1_65___stage___block_26_v_x = _q___pip_5160_1_65___stage___block_26_v_x;
_d___pip_5160_1_66___stage___block_26_v_x = _q___pip_5160_1_66___stage___block_26_v_x;
_d___pip_5160_1_67___stage___block_26_v_x = _q___pip_5160_1_67___stage___block_26_v_x;
_d___pip_5160_1_68___stage___block_26_v_x = _q___pip_5160_1_68___stage___block_26_v_x;
_d___pip_5160_1_69___stage___block_26_v_x = _q___pip_5160_1_69___stage___block_26_v_x;
_d___pip_5160_1_70___stage___block_26_v_x = _q___pip_5160_1_70___stage___block_26_v_x;
_d___pip_5160_1_71___stage___block_26_v_x = _q___pip_5160_1_71___stage___block_26_v_x;
_d___pip_5160_1_72___stage___block_26_v_x = _q___pip_5160_1_72___stage___block_26_v_x;
_d___pip_5160_1_73___stage___block_26_v_x = _q___pip_5160_1_73___stage___block_26_v_x;
_d___pip_5160_1_74___stage___block_26_v_x = _q___pip_5160_1_74___stage___block_26_v_x;
_d___pip_5160_1_75___stage___block_26_v_x = _q___pip_5160_1_75___stage___block_26_v_x;
_d___pip_5160_1_76___stage___block_26_v_x = _q___pip_5160_1_76___stage___block_26_v_x;
_d___pip_5160_1_77___stage___block_26_v_x = _q___pip_5160_1_77___stage___block_26_v_x;
_d___pip_5160_1_78___stage___block_26_v_x = _q___pip_5160_1_78___stage___block_26_v_x;
_d___pip_5160_1_79___stage___block_26_v_x = _q___pip_5160_1_79___stage___block_26_v_x;
_d___pip_5160_1_80___stage___block_26_v_x = _q___pip_5160_1_80___stage___block_26_v_x;
_d___pip_5160_1_81___stage___block_26_v_x = _q___pip_5160_1_81___stage___block_26_v_x;
_d___pip_5160_1_82___stage___block_26_v_x = _q___pip_5160_1_82___stage___block_26_v_x;
_d___pip_5160_1_83___stage___block_26_v_x = _q___pip_5160_1_83___stage___block_26_v_x;
_d___pip_5160_1_84___stage___block_26_v_x = _q___pip_5160_1_84___stage___block_26_v_x;
_d___pip_5160_1_85___stage___block_26_v_x = _q___pip_5160_1_85___stage___block_26_v_x;
_d___pip_5160_1_86___stage___block_26_v_x = _q___pip_5160_1_86___stage___block_26_v_x;
_d___pip_5160_1_87___stage___block_26_v_x = _q___pip_5160_1_87___stage___block_26_v_x;
_d___pip_5160_1_88___stage___block_26_v_x = _q___pip_5160_1_88___stage___block_26_v_x;
_d___pip_5160_1_89___stage___block_26_v_x = _q___pip_5160_1_89___stage___block_26_v_x;
_d___pip_5160_1_90___stage___block_26_v_x = _q___pip_5160_1_90___stage___block_26_v_x;
_d___pip_5160_1_91___stage___block_26_v_x = _q___pip_5160_1_91___stage___block_26_v_x;
_d___pip_5160_1_92___stage___block_26_v_x = _q___pip_5160_1_92___stage___block_26_v_x;
_d___pip_5160_1_93___stage___block_26_v_x = _q___pip_5160_1_93___stage___block_26_v_x;
_d___pip_5160_1_94___stage___block_26_v_x = _q___pip_5160_1_94___stage___block_26_v_x;
_d___pip_5160_1_95___stage___block_26_v_x = _q___pip_5160_1_95___stage___block_26_v_x;
_d___pip_5160_1_96___stage___block_26_v_x = _q___pip_5160_1_96___stage___block_26_v_x;
_d___pip_5160_1_97___stage___block_26_v_x = _q___pip_5160_1_97___stage___block_26_v_x;
_d___pip_5160_1_98___stage___block_26_v_x = _q___pip_5160_1_98___stage___block_26_v_x;
_d___pip_5160_1_99___stage___block_26_v_x = _q___pip_5160_1_99___stage___block_26_v_x;
_d___pip_5160_1_100___stage___block_26_v_x = _q___pip_5160_1_100___stage___block_26_v_x;
_d___pip_5160_1_101___stage___block_26_v_x = _q___pip_5160_1_101___stage___block_26_v_x;
_d___pip_5160_1_102___stage___block_26_v_x = _q___pip_5160_1_102___stage___block_26_v_x;
_d___pip_5160_1_103___stage___block_26_v_x = _q___pip_5160_1_103___stage___block_26_v_x;
_d___pip_5160_1_104___stage___block_26_v_x = _q___pip_5160_1_104___stage___block_26_v_x;
_d___pip_5160_1_105___stage___block_26_v_x = _q___pip_5160_1_105___stage___block_26_v_x;
_d___pip_5160_1_106___stage___block_26_v_x = _q___pip_5160_1_106___stage___block_26_v_x;
_d___pip_5160_1_107___stage___block_26_v_x = _q___pip_5160_1_107___stage___block_26_v_x;
_d___pip_5160_1_108___stage___block_26_v_x = _q___pip_5160_1_108___stage___block_26_v_x;
_d___pip_5160_1_109___stage___block_26_v_x = _q___pip_5160_1_109___stage___block_26_v_x;
_d___pip_5160_1_110___stage___block_26_v_x = _q___pip_5160_1_110___stage___block_26_v_x;
_d___pip_5160_1_111___stage___block_26_v_x = _q___pip_5160_1_111___stage___block_26_v_x;
_d___pip_5160_1_112___stage___block_26_v_x = _q___pip_5160_1_112___stage___block_26_v_x;
_d___pip_5160_1_113___stage___block_26_v_x = _q___pip_5160_1_113___stage___block_26_v_x;
_d___pip_5160_1_114___stage___block_26_v_x = _q___pip_5160_1_114___stage___block_26_v_x;
_d___pip_5160_1_115___stage___block_26_v_x = _q___pip_5160_1_115___stage___block_26_v_x;
_d___pip_5160_1_116___stage___block_26_v_x = _q___pip_5160_1_116___stage___block_26_v_x;
_d___pip_5160_1_117___stage___block_26_v_x = _q___pip_5160_1_117___stage___block_26_v_x;
_d___pip_5160_1_118___stage___block_26_v_x = _q___pip_5160_1_118___stage___block_26_v_x;
_d___pip_5160_1_119___stage___block_26_v_x = _q___pip_5160_1_119___stage___block_26_v_x;
_d___pip_5160_1_120___stage___block_26_v_x = _q___pip_5160_1_120___stage___block_26_v_x;
_d___pip_5160_1_121___stage___block_26_v_x = _q___pip_5160_1_121___stage___block_26_v_x;
_d___pip_5160_1_122___stage___block_26_v_x = _q___pip_5160_1_122___stage___block_26_v_x;
_d___pip_5160_1_123___stage___block_26_v_x = _q___pip_5160_1_123___stage___block_26_v_x;
_d___pip_5160_1_124___stage___block_26_v_x = _q___pip_5160_1_124___stage___block_26_v_x;
_d___pip_5160_1_125___stage___block_26_v_x = _q___pip_5160_1_125___stage___block_26_v_x;
_d___pip_5160_1_126___stage___block_26_v_x = _q___pip_5160_1_126___stage___block_26_v_x;
_d___pip_5160_1_127___stage___block_26_v_x = _q___pip_5160_1_127___stage___block_26_v_x;
_d___pip_5160_1_128___stage___block_26_v_x = _q___pip_5160_1_128___stage___block_26_v_x;
_d___pip_5160_1_129___stage___block_26_v_x = _q___pip_5160_1_129___stage___block_26_v_x;
_d___pip_5160_1_130___stage___block_26_v_x = _q___pip_5160_1_130___stage___block_26_v_x;
_d___pip_5160_1_131___stage___block_26_v_x = _q___pip_5160_1_131___stage___block_26_v_x;
_d___pip_5160_1_132___stage___block_26_v_x = _q___pip_5160_1_132___stage___block_26_v_x;
_d___pip_5160_1_133___stage___block_26_v_x = _q___pip_5160_1_133___stage___block_26_v_x;
_d___pip_5160_1_134___stage___block_26_v_x = _q___pip_5160_1_134___stage___block_26_v_x;
_d___pip_5160_1_4___stage___block_26_v_y = _q___pip_5160_1_4___stage___block_26_v_y;
_d___pip_5160_1_5___stage___block_26_v_y = _q___pip_5160_1_5___stage___block_26_v_y;
_d___pip_5160_1_6___stage___block_26_v_y = _q___pip_5160_1_6___stage___block_26_v_y;
_d___pip_5160_1_7___stage___block_26_v_y = _q___pip_5160_1_7___stage___block_26_v_y;
_d___pip_5160_1_8___stage___block_26_v_y = _q___pip_5160_1_8___stage___block_26_v_y;
_d___pip_5160_1_9___stage___block_26_v_y = _q___pip_5160_1_9___stage___block_26_v_y;
_d___pip_5160_1_10___stage___block_26_v_y = _q___pip_5160_1_10___stage___block_26_v_y;
_d___pip_5160_1_11___stage___block_26_v_y = _q___pip_5160_1_11___stage___block_26_v_y;
_d___pip_5160_1_12___stage___block_26_v_y = _q___pip_5160_1_12___stage___block_26_v_y;
_d___pip_5160_1_13___stage___block_26_v_y = _q___pip_5160_1_13___stage___block_26_v_y;
_d___pip_5160_1_14___stage___block_26_v_y = _q___pip_5160_1_14___stage___block_26_v_y;
_d___pip_5160_1_15___stage___block_26_v_y = _q___pip_5160_1_15___stage___block_26_v_y;
_d___pip_5160_1_16___stage___block_26_v_y = _q___pip_5160_1_16___stage___block_26_v_y;
_d___pip_5160_1_17___stage___block_26_v_y = _q___pip_5160_1_17___stage___block_26_v_y;
_d___pip_5160_1_18___stage___block_26_v_y = _q___pip_5160_1_18___stage___block_26_v_y;
_d___pip_5160_1_19___stage___block_26_v_y = _q___pip_5160_1_19___stage___block_26_v_y;
_d___pip_5160_1_20___stage___block_26_v_y = _q___pip_5160_1_20___stage___block_26_v_y;
_d___pip_5160_1_21___stage___block_26_v_y = _q___pip_5160_1_21___stage___block_26_v_y;
_d___pip_5160_1_22___stage___block_26_v_y = _q___pip_5160_1_22___stage___block_26_v_y;
_d___pip_5160_1_23___stage___block_26_v_y = _q___pip_5160_1_23___stage___block_26_v_y;
_d___pip_5160_1_24___stage___block_26_v_y = _q___pip_5160_1_24___stage___block_26_v_y;
_d___pip_5160_1_25___stage___block_26_v_y = _q___pip_5160_1_25___stage___block_26_v_y;
_d___pip_5160_1_26___stage___block_26_v_y = _q___pip_5160_1_26___stage___block_26_v_y;
_d___pip_5160_1_27___stage___block_26_v_y = _q___pip_5160_1_27___stage___block_26_v_y;
_d___pip_5160_1_28___stage___block_26_v_y = _q___pip_5160_1_28___stage___block_26_v_y;
_d___pip_5160_1_29___stage___block_26_v_y = _q___pip_5160_1_29___stage___block_26_v_y;
_d___pip_5160_1_30___stage___block_26_v_y = _q___pip_5160_1_30___stage___block_26_v_y;
_d___pip_5160_1_31___stage___block_26_v_y = _q___pip_5160_1_31___stage___block_26_v_y;
_d___pip_5160_1_32___stage___block_26_v_y = _q___pip_5160_1_32___stage___block_26_v_y;
_d___pip_5160_1_33___stage___block_26_v_y = _q___pip_5160_1_33___stage___block_26_v_y;
_d___pip_5160_1_34___stage___block_26_v_y = _q___pip_5160_1_34___stage___block_26_v_y;
_d___pip_5160_1_35___stage___block_26_v_y = _q___pip_5160_1_35___stage___block_26_v_y;
_d___pip_5160_1_36___stage___block_26_v_y = _q___pip_5160_1_36___stage___block_26_v_y;
_d___pip_5160_1_37___stage___block_26_v_y = _q___pip_5160_1_37___stage___block_26_v_y;
_d___pip_5160_1_38___stage___block_26_v_y = _q___pip_5160_1_38___stage___block_26_v_y;
_d___pip_5160_1_39___stage___block_26_v_y = _q___pip_5160_1_39___stage___block_26_v_y;
_d___pip_5160_1_40___stage___block_26_v_y = _q___pip_5160_1_40___stage___block_26_v_y;
_d___pip_5160_1_41___stage___block_26_v_y = _q___pip_5160_1_41___stage___block_26_v_y;
_d___pip_5160_1_42___stage___block_26_v_y = _q___pip_5160_1_42___stage___block_26_v_y;
_d___pip_5160_1_43___stage___block_26_v_y = _q___pip_5160_1_43___stage___block_26_v_y;
_d___pip_5160_1_44___stage___block_26_v_y = _q___pip_5160_1_44___stage___block_26_v_y;
_d___pip_5160_1_45___stage___block_26_v_y = _q___pip_5160_1_45___stage___block_26_v_y;
_d___pip_5160_1_46___stage___block_26_v_y = _q___pip_5160_1_46___stage___block_26_v_y;
_d___pip_5160_1_47___stage___block_26_v_y = _q___pip_5160_1_47___stage___block_26_v_y;
_d___pip_5160_1_48___stage___block_26_v_y = _q___pip_5160_1_48___stage___block_26_v_y;
_d___pip_5160_1_49___stage___block_26_v_y = _q___pip_5160_1_49___stage___block_26_v_y;
_d___pip_5160_1_50___stage___block_26_v_y = _q___pip_5160_1_50___stage___block_26_v_y;
_d___pip_5160_1_51___stage___block_26_v_y = _q___pip_5160_1_51___stage___block_26_v_y;
_d___pip_5160_1_52___stage___block_26_v_y = _q___pip_5160_1_52___stage___block_26_v_y;
_d___pip_5160_1_53___stage___block_26_v_y = _q___pip_5160_1_53___stage___block_26_v_y;
_d___pip_5160_1_54___stage___block_26_v_y = _q___pip_5160_1_54___stage___block_26_v_y;
_d___pip_5160_1_55___stage___block_26_v_y = _q___pip_5160_1_55___stage___block_26_v_y;
_d___pip_5160_1_56___stage___block_26_v_y = _q___pip_5160_1_56___stage___block_26_v_y;
_d___pip_5160_1_57___stage___block_26_v_y = _q___pip_5160_1_57___stage___block_26_v_y;
_d___pip_5160_1_58___stage___block_26_v_y = _q___pip_5160_1_58___stage___block_26_v_y;
_d___pip_5160_1_59___stage___block_26_v_y = _q___pip_5160_1_59___stage___block_26_v_y;
_d___pip_5160_1_60___stage___block_26_v_y = _q___pip_5160_1_60___stage___block_26_v_y;
_d___pip_5160_1_61___stage___block_26_v_y = _q___pip_5160_1_61___stage___block_26_v_y;
_d___pip_5160_1_62___stage___block_26_v_y = _q___pip_5160_1_62___stage___block_26_v_y;
_d___pip_5160_1_63___stage___block_26_v_y = _q___pip_5160_1_63___stage___block_26_v_y;
_d___pip_5160_1_64___stage___block_26_v_y = _q___pip_5160_1_64___stage___block_26_v_y;
_d___pip_5160_1_65___stage___block_26_v_y = _q___pip_5160_1_65___stage___block_26_v_y;
_d___pip_5160_1_66___stage___block_26_v_y = _q___pip_5160_1_66___stage___block_26_v_y;
_d___pip_5160_1_67___stage___block_26_v_y = _q___pip_5160_1_67___stage___block_26_v_y;
_d___pip_5160_1_68___stage___block_26_v_y = _q___pip_5160_1_68___stage___block_26_v_y;
_d___pip_5160_1_69___stage___block_26_v_y = _q___pip_5160_1_69___stage___block_26_v_y;
_d___pip_5160_1_70___stage___block_26_v_y = _q___pip_5160_1_70___stage___block_26_v_y;
_d___pip_5160_1_71___stage___block_26_v_y = _q___pip_5160_1_71___stage___block_26_v_y;
_d___pip_5160_1_72___stage___block_26_v_y = _q___pip_5160_1_72___stage___block_26_v_y;
_d___pip_5160_1_73___stage___block_26_v_y = _q___pip_5160_1_73___stage___block_26_v_y;
_d___pip_5160_1_74___stage___block_26_v_y = _q___pip_5160_1_74___stage___block_26_v_y;
_d___pip_5160_1_75___stage___block_26_v_y = _q___pip_5160_1_75___stage___block_26_v_y;
_d___pip_5160_1_76___stage___block_26_v_y = _q___pip_5160_1_76___stage___block_26_v_y;
_d___pip_5160_1_77___stage___block_26_v_y = _q___pip_5160_1_77___stage___block_26_v_y;
_d___pip_5160_1_78___stage___block_26_v_y = _q___pip_5160_1_78___stage___block_26_v_y;
_d___pip_5160_1_79___stage___block_26_v_y = _q___pip_5160_1_79___stage___block_26_v_y;
_d___pip_5160_1_80___stage___block_26_v_y = _q___pip_5160_1_80___stage___block_26_v_y;
_d___pip_5160_1_81___stage___block_26_v_y = _q___pip_5160_1_81___stage___block_26_v_y;
_d___pip_5160_1_82___stage___block_26_v_y = _q___pip_5160_1_82___stage___block_26_v_y;
_d___pip_5160_1_83___stage___block_26_v_y = _q___pip_5160_1_83___stage___block_26_v_y;
_d___pip_5160_1_84___stage___block_26_v_y = _q___pip_5160_1_84___stage___block_26_v_y;
_d___pip_5160_1_85___stage___block_26_v_y = _q___pip_5160_1_85___stage___block_26_v_y;
_d___pip_5160_1_86___stage___block_26_v_y = _q___pip_5160_1_86___stage___block_26_v_y;
_d___pip_5160_1_87___stage___block_26_v_y = _q___pip_5160_1_87___stage___block_26_v_y;
_d___pip_5160_1_88___stage___block_26_v_y = _q___pip_5160_1_88___stage___block_26_v_y;
_d___pip_5160_1_89___stage___block_26_v_y = _q___pip_5160_1_89___stage___block_26_v_y;
_d___pip_5160_1_90___stage___block_26_v_y = _q___pip_5160_1_90___stage___block_26_v_y;
_d___pip_5160_1_91___stage___block_26_v_y = _q___pip_5160_1_91___stage___block_26_v_y;
_d___pip_5160_1_92___stage___block_26_v_y = _q___pip_5160_1_92___stage___block_26_v_y;
_d___pip_5160_1_93___stage___block_26_v_y = _q___pip_5160_1_93___stage___block_26_v_y;
_d___pip_5160_1_94___stage___block_26_v_y = _q___pip_5160_1_94___stage___block_26_v_y;
_d___pip_5160_1_95___stage___block_26_v_y = _q___pip_5160_1_95___stage___block_26_v_y;
_d___pip_5160_1_96___stage___block_26_v_y = _q___pip_5160_1_96___stage___block_26_v_y;
_d___pip_5160_1_97___stage___block_26_v_y = _q___pip_5160_1_97___stage___block_26_v_y;
_d___pip_5160_1_98___stage___block_26_v_y = _q___pip_5160_1_98___stage___block_26_v_y;
_d___pip_5160_1_99___stage___block_26_v_y = _q___pip_5160_1_99___stage___block_26_v_y;
_d___pip_5160_1_100___stage___block_26_v_y = _q___pip_5160_1_100___stage___block_26_v_y;
_d___pip_5160_1_101___stage___block_26_v_y = _q___pip_5160_1_101___stage___block_26_v_y;
_d___pip_5160_1_102___stage___block_26_v_y = _q___pip_5160_1_102___stage___block_26_v_y;
_d___pip_5160_1_103___stage___block_26_v_y = _q___pip_5160_1_103___stage___block_26_v_y;
_d___pip_5160_1_104___stage___block_26_v_y = _q___pip_5160_1_104___stage___block_26_v_y;
_d___pip_5160_1_105___stage___block_26_v_y = _q___pip_5160_1_105___stage___block_26_v_y;
_d___pip_5160_1_106___stage___block_26_v_y = _q___pip_5160_1_106___stage___block_26_v_y;
_d___pip_5160_1_107___stage___block_26_v_y = _q___pip_5160_1_107___stage___block_26_v_y;
_d___pip_5160_1_108___stage___block_26_v_y = _q___pip_5160_1_108___stage___block_26_v_y;
_d___pip_5160_1_109___stage___block_26_v_y = _q___pip_5160_1_109___stage___block_26_v_y;
_d___pip_5160_1_110___stage___block_26_v_y = _q___pip_5160_1_110___stage___block_26_v_y;
_d___pip_5160_1_111___stage___block_26_v_y = _q___pip_5160_1_111___stage___block_26_v_y;
_d___pip_5160_1_112___stage___block_26_v_y = _q___pip_5160_1_112___stage___block_26_v_y;
_d___pip_5160_1_113___stage___block_26_v_y = _q___pip_5160_1_113___stage___block_26_v_y;
_d___pip_5160_1_114___stage___block_26_v_y = _q___pip_5160_1_114___stage___block_26_v_y;
_d___pip_5160_1_115___stage___block_26_v_y = _q___pip_5160_1_115___stage___block_26_v_y;
_d___pip_5160_1_116___stage___block_26_v_y = _q___pip_5160_1_116___stage___block_26_v_y;
_d___pip_5160_1_117___stage___block_26_v_y = _q___pip_5160_1_117___stage___block_26_v_y;
_d___pip_5160_1_118___stage___block_26_v_y = _q___pip_5160_1_118___stage___block_26_v_y;
_d___pip_5160_1_119___stage___block_26_v_y = _q___pip_5160_1_119___stage___block_26_v_y;
_d___pip_5160_1_120___stage___block_26_v_y = _q___pip_5160_1_120___stage___block_26_v_y;
_d___pip_5160_1_121___stage___block_26_v_y = _q___pip_5160_1_121___stage___block_26_v_y;
_d___pip_5160_1_122___stage___block_26_v_y = _q___pip_5160_1_122___stage___block_26_v_y;
_d___pip_5160_1_123___stage___block_26_v_y = _q___pip_5160_1_123___stage___block_26_v_y;
_d___pip_5160_1_124___stage___block_26_v_y = _q___pip_5160_1_124___stage___block_26_v_y;
_d___pip_5160_1_125___stage___block_26_v_y = _q___pip_5160_1_125___stage___block_26_v_y;
_d___pip_5160_1_126___stage___block_26_v_y = _q___pip_5160_1_126___stage___block_26_v_y;
_d___pip_5160_1_127___stage___block_26_v_y = _q___pip_5160_1_127___stage___block_26_v_y;
_d___pip_5160_1_128___stage___block_26_v_y = _q___pip_5160_1_128___stage___block_26_v_y;
_d___pip_5160_1_129___stage___block_26_v_y = _q___pip_5160_1_129___stage___block_26_v_y;
_d___pip_5160_1_130___stage___block_26_v_y = _q___pip_5160_1_130___stage___block_26_v_y;
_d___pip_5160_1_131___stage___block_26_v_y = _q___pip_5160_1_131___stage___block_26_v_y;
_d___pip_5160_1_132___stage___block_26_v_y = _q___pip_5160_1_132___stage___block_26_v_y;
_d___pip_5160_1_133___stage___block_26_v_y = _q___pip_5160_1_133___stage___block_26_v_y;
_d___pip_5160_1_134___stage___block_26_v_y = _q___pip_5160_1_134___stage___block_26_v_y;
_d___pip_5160_1_4___stage___block_26_v_z = _q___pip_5160_1_4___stage___block_26_v_z;
_d___pip_5160_1_5___stage___block_26_v_z = _q___pip_5160_1_5___stage___block_26_v_z;
_d___pip_5160_1_6___stage___block_26_v_z = _q___pip_5160_1_6___stage___block_26_v_z;
_d___pip_5160_1_7___stage___block_26_v_z = _q___pip_5160_1_7___stage___block_26_v_z;
_d___pip_5160_1_8___stage___block_26_v_z = _q___pip_5160_1_8___stage___block_26_v_z;
_d___pip_5160_1_9___stage___block_26_v_z = _q___pip_5160_1_9___stage___block_26_v_z;
_d___pip_5160_1_10___stage___block_26_v_z = _q___pip_5160_1_10___stage___block_26_v_z;
_d___pip_5160_1_11___stage___block_26_v_z = _q___pip_5160_1_11___stage___block_26_v_z;
_d___pip_5160_1_12___stage___block_26_v_z = _q___pip_5160_1_12___stage___block_26_v_z;
_d___pip_5160_1_13___stage___block_26_v_z = _q___pip_5160_1_13___stage___block_26_v_z;
_d___pip_5160_1_14___stage___block_26_v_z = _q___pip_5160_1_14___stage___block_26_v_z;
_d___pip_5160_1_15___stage___block_26_v_z = _q___pip_5160_1_15___stage___block_26_v_z;
_d___pip_5160_1_16___stage___block_26_v_z = _q___pip_5160_1_16___stage___block_26_v_z;
_d___pip_5160_1_17___stage___block_26_v_z = _q___pip_5160_1_17___stage___block_26_v_z;
_d___pip_5160_1_18___stage___block_26_v_z = _q___pip_5160_1_18___stage___block_26_v_z;
_d___pip_5160_1_19___stage___block_26_v_z = _q___pip_5160_1_19___stage___block_26_v_z;
_d___pip_5160_1_20___stage___block_26_v_z = _q___pip_5160_1_20___stage___block_26_v_z;
_d___pip_5160_1_21___stage___block_26_v_z = _q___pip_5160_1_21___stage___block_26_v_z;
_d___pip_5160_1_22___stage___block_26_v_z = _q___pip_5160_1_22___stage___block_26_v_z;
_d___pip_5160_1_23___stage___block_26_v_z = _q___pip_5160_1_23___stage___block_26_v_z;
_d___pip_5160_1_24___stage___block_26_v_z = _q___pip_5160_1_24___stage___block_26_v_z;
_d___pip_5160_1_25___stage___block_26_v_z = _q___pip_5160_1_25___stage___block_26_v_z;
_d___pip_5160_1_26___stage___block_26_v_z = _q___pip_5160_1_26___stage___block_26_v_z;
_d___pip_5160_1_27___stage___block_26_v_z = _q___pip_5160_1_27___stage___block_26_v_z;
_d___pip_5160_1_28___stage___block_26_v_z = _q___pip_5160_1_28___stage___block_26_v_z;
_d___pip_5160_1_29___stage___block_26_v_z = _q___pip_5160_1_29___stage___block_26_v_z;
_d___pip_5160_1_30___stage___block_26_v_z = _q___pip_5160_1_30___stage___block_26_v_z;
_d___pip_5160_1_31___stage___block_26_v_z = _q___pip_5160_1_31___stage___block_26_v_z;
_d___pip_5160_1_32___stage___block_26_v_z = _q___pip_5160_1_32___stage___block_26_v_z;
_d___pip_5160_1_33___stage___block_26_v_z = _q___pip_5160_1_33___stage___block_26_v_z;
_d___pip_5160_1_34___stage___block_26_v_z = _q___pip_5160_1_34___stage___block_26_v_z;
_d___pip_5160_1_35___stage___block_26_v_z = _q___pip_5160_1_35___stage___block_26_v_z;
_d___pip_5160_1_36___stage___block_26_v_z = _q___pip_5160_1_36___stage___block_26_v_z;
_d___pip_5160_1_37___stage___block_26_v_z = _q___pip_5160_1_37___stage___block_26_v_z;
_d___pip_5160_1_38___stage___block_26_v_z = _q___pip_5160_1_38___stage___block_26_v_z;
_d___pip_5160_1_39___stage___block_26_v_z = _q___pip_5160_1_39___stage___block_26_v_z;
_d___pip_5160_1_40___stage___block_26_v_z = _q___pip_5160_1_40___stage___block_26_v_z;
_d___pip_5160_1_41___stage___block_26_v_z = _q___pip_5160_1_41___stage___block_26_v_z;
_d___pip_5160_1_42___stage___block_26_v_z = _q___pip_5160_1_42___stage___block_26_v_z;
_d___pip_5160_1_43___stage___block_26_v_z = _q___pip_5160_1_43___stage___block_26_v_z;
_d___pip_5160_1_44___stage___block_26_v_z = _q___pip_5160_1_44___stage___block_26_v_z;
_d___pip_5160_1_45___stage___block_26_v_z = _q___pip_5160_1_45___stage___block_26_v_z;
_d___pip_5160_1_46___stage___block_26_v_z = _q___pip_5160_1_46___stage___block_26_v_z;
_d___pip_5160_1_47___stage___block_26_v_z = _q___pip_5160_1_47___stage___block_26_v_z;
_d___pip_5160_1_48___stage___block_26_v_z = _q___pip_5160_1_48___stage___block_26_v_z;
_d___pip_5160_1_49___stage___block_26_v_z = _q___pip_5160_1_49___stage___block_26_v_z;
_d___pip_5160_1_50___stage___block_26_v_z = _q___pip_5160_1_50___stage___block_26_v_z;
_d___pip_5160_1_51___stage___block_26_v_z = _q___pip_5160_1_51___stage___block_26_v_z;
_d___pip_5160_1_52___stage___block_26_v_z = _q___pip_5160_1_52___stage___block_26_v_z;
_d___pip_5160_1_53___stage___block_26_v_z = _q___pip_5160_1_53___stage___block_26_v_z;
_d___pip_5160_1_54___stage___block_26_v_z = _q___pip_5160_1_54___stage___block_26_v_z;
_d___pip_5160_1_55___stage___block_26_v_z = _q___pip_5160_1_55___stage___block_26_v_z;
_d___pip_5160_1_56___stage___block_26_v_z = _q___pip_5160_1_56___stage___block_26_v_z;
_d___pip_5160_1_57___stage___block_26_v_z = _q___pip_5160_1_57___stage___block_26_v_z;
_d___pip_5160_1_58___stage___block_26_v_z = _q___pip_5160_1_58___stage___block_26_v_z;
_d___pip_5160_1_59___stage___block_26_v_z = _q___pip_5160_1_59___stage___block_26_v_z;
_d___pip_5160_1_60___stage___block_26_v_z = _q___pip_5160_1_60___stage___block_26_v_z;
_d___pip_5160_1_61___stage___block_26_v_z = _q___pip_5160_1_61___stage___block_26_v_z;
_d___pip_5160_1_62___stage___block_26_v_z = _q___pip_5160_1_62___stage___block_26_v_z;
_d___pip_5160_1_63___stage___block_26_v_z = _q___pip_5160_1_63___stage___block_26_v_z;
_d___pip_5160_1_64___stage___block_26_v_z = _q___pip_5160_1_64___stage___block_26_v_z;
_d___pip_5160_1_65___stage___block_26_v_z = _q___pip_5160_1_65___stage___block_26_v_z;
_d___pip_5160_1_66___stage___block_26_v_z = _q___pip_5160_1_66___stage___block_26_v_z;
_d___pip_5160_1_67___stage___block_26_v_z = _q___pip_5160_1_67___stage___block_26_v_z;
_d___pip_5160_1_68___stage___block_26_v_z = _q___pip_5160_1_68___stage___block_26_v_z;
_d___pip_5160_1_69___stage___block_26_v_z = _q___pip_5160_1_69___stage___block_26_v_z;
_d___pip_5160_1_70___stage___block_26_v_z = _q___pip_5160_1_70___stage___block_26_v_z;
_d___pip_5160_1_71___stage___block_26_v_z = _q___pip_5160_1_71___stage___block_26_v_z;
_d___pip_5160_1_72___stage___block_26_v_z = _q___pip_5160_1_72___stage___block_26_v_z;
_d___pip_5160_1_73___stage___block_26_v_z = _q___pip_5160_1_73___stage___block_26_v_z;
_d___pip_5160_1_74___stage___block_26_v_z = _q___pip_5160_1_74___stage___block_26_v_z;
_d___pip_5160_1_75___stage___block_26_v_z = _q___pip_5160_1_75___stage___block_26_v_z;
_d___pip_5160_1_76___stage___block_26_v_z = _q___pip_5160_1_76___stage___block_26_v_z;
_d___pip_5160_1_77___stage___block_26_v_z = _q___pip_5160_1_77___stage___block_26_v_z;
_d___pip_5160_1_78___stage___block_26_v_z = _q___pip_5160_1_78___stage___block_26_v_z;
_d___pip_5160_1_79___stage___block_26_v_z = _q___pip_5160_1_79___stage___block_26_v_z;
_d___pip_5160_1_80___stage___block_26_v_z = _q___pip_5160_1_80___stage___block_26_v_z;
_d___pip_5160_1_81___stage___block_26_v_z = _q___pip_5160_1_81___stage___block_26_v_z;
_d___pip_5160_1_82___stage___block_26_v_z = _q___pip_5160_1_82___stage___block_26_v_z;
_d___pip_5160_1_83___stage___block_26_v_z = _q___pip_5160_1_83___stage___block_26_v_z;
_d___pip_5160_1_84___stage___block_26_v_z = _q___pip_5160_1_84___stage___block_26_v_z;
_d___pip_5160_1_85___stage___block_26_v_z = _q___pip_5160_1_85___stage___block_26_v_z;
_d___pip_5160_1_86___stage___block_26_v_z = _q___pip_5160_1_86___stage___block_26_v_z;
_d___pip_5160_1_87___stage___block_26_v_z = _q___pip_5160_1_87___stage___block_26_v_z;
_d___pip_5160_1_88___stage___block_26_v_z = _q___pip_5160_1_88___stage___block_26_v_z;
_d___pip_5160_1_89___stage___block_26_v_z = _q___pip_5160_1_89___stage___block_26_v_z;
_d___pip_5160_1_90___stage___block_26_v_z = _q___pip_5160_1_90___stage___block_26_v_z;
_d___pip_5160_1_91___stage___block_26_v_z = _q___pip_5160_1_91___stage___block_26_v_z;
_d___pip_5160_1_92___stage___block_26_v_z = _q___pip_5160_1_92___stage___block_26_v_z;
_d___pip_5160_1_93___stage___block_26_v_z = _q___pip_5160_1_93___stage___block_26_v_z;
_d___pip_5160_1_94___stage___block_26_v_z = _q___pip_5160_1_94___stage___block_26_v_z;
_d___pip_5160_1_95___stage___block_26_v_z = _q___pip_5160_1_95___stage___block_26_v_z;
_d___pip_5160_1_96___stage___block_26_v_z = _q___pip_5160_1_96___stage___block_26_v_z;
_d___pip_5160_1_97___stage___block_26_v_z = _q___pip_5160_1_97___stage___block_26_v_z;
_d___pip_5160_1_98___stage___block_26_v_z = _q___pip_5160_1_98___stage___block_26_v_z;
_d___pip_5160_1_99___stage___block_26_v_z = _q___pip_5160_1_99___stage___block_26_v_z;
_d___pip_5160_1_100___stage___block_26_v_z = _q___pip_5160_1_100___stage___block_26_v_z;
_d___pip_5160_1_101___stage___block_26_v_z = _q___pip_5160_1_101___stage___block_26_v_z;
_d___pip_5160_1_102___stage___block_26_v_z = _q___pip_5160_1_102___stage___block_26_v_z;
_d___pip_5160_1_103___stage___block_26_v_z = _q___pip_5160_1_103___stage___block_26_v_z;
_d___pip_5160_1_104___stage___block_26_v_z = _q___pip_5160_1_104___stage___block_26_v_z;
_d___pip_5160_1_105___stage___block_26_v_z = _q___pip_5160_1_105___stage___block_26_v_z;
_d___pip_5160_1_106___stage___block_26_v_z = _q___pip_5160_1_106___stage___block_26_v_z;
_d___pip_5160_1_107___stage___block_26_v_z = _q___pip_5160_1_107___stage___block_26_v_z;
_d___pip_5160_1_108___stage___block_26_v_z = _q___pip_5160_1_108___stage___block_26_v_z;
_d___pip_5160_1_109___stage___block_26_v_z = _q___pip_5160_1_109___stage___block_26_v_z;
_d___pip_5160_1_110___stage___block_26_v_z = _q___pip_5160_1_110___stage___block_26_v_z;
_d___pip_5160_1_111___stage___block_26_v_z = _q___pip_5160_1_111___stage___block_26_v_z;
_d___pip_5160_1_112___stage___block_26_v_z = _q___pip_5160_1_112___stage___block_26_v_z;
_d___pip_5160_1_113___stage___block_26_v_z = _q___pip_5160_1_113___stage___block_26_v_z;
_d___pip_5160_1_114___stage___block_26_v_z = _q___pip_5160_1_114___stage___block_26_v_z;
_d___pip_5160_1_115___stage___block_26_v_z = _q___pip_5160_1_115___stage___block_26_v_z;
_d___pip_5160_1_116___stage___block_26_v_z = _q___pip_5160_1_116___stage___block_26_v_z;
_d___pip_5160_1_117___stage___block_26_v_z = _q___pip_5160_1_117___stage___block_26_v_z;
_d___pip_5160_1_118___stage___block_26_v_z = _q___pip_5160_1_118___stage___block_26_v_z;
_d___pip_5160_1_119___stage___block_26_v_z = _q___pip_5160_1_119___stage___block_26_v_z;
_d___pip_5160_1_120___stage___block_26_v_z = _q___pip_5160_1_120___stage___block_26_v_z;
_d___pip_5160_1_121___stage___block_26_v_z = _q___pip_5160_1_121___stage___block_26_v_z;
_d___pip_5160_1_122___stage___block_26_v_z = _q___pip_5160_1_122___stage___block_26_v_z;
_d___pip_5160_1_123___stage___block_26_v_z = _q___pip_5160_1_123___stage___block_26_v_z;
_d___pip_5160_1_124___stage___block_26_v_z = _q___pip_5160_1_124___stage___block_26_v_z;
_d___pip_5160_1_125___stage___block_26_v_z = _q___pip_5160_1_125___stage___block_26_v_z;
_d___pip_5160_1_126___stage___block_26_v_z = _q___pip_5160_1_126___stage___block_26_v_z;
_d___pip_5160_1_127___stage___block_26_v_z = _q___pip_5160_1_127___stage___block_26_v_z;
_d___pip_5160_1_128___stage___block_26_v_z = _q___pip_5160_1_128___stage___block_26_v_z;
_d___pip_5160_1_129___stage___block_26_v_z = _q___pip_5160_1_129___stage___block_26_v_z;
_d___pip_5160_1_130___stage___block_26_v_z = _q___pip_5160_1_130___stage___block_26_v_z;
_d___pip_5160_1_131___stage___block_26_v_z = _q___pip_5160_1_131___stage___block_26_v_z;
_d___pip_5160_1_132___stage___block_26_v_z = _q___pip_5160_1_132___stage___block_26_v_z;
_d___pip_5160_1_133___stage___block_26_v_z = _q___pip_5160_1_133___stage___block_26_v_z;
_d___pip_5160_1_134___stage___block_26_v_z = _q___pip_5160_1_134___stage___block_26_v_z;
_d___pip_5160_1_0___stage___block_6_clr = _q___pip_5160_1_0___stage___block_6_clr;
_d___pip_5160_1_1___stage___block_6_clr = _q___pip_5160_1_1___stage___block_6_clr;
_d___pip_5160_1_2___stage___block_6_clr = _q___pip_5160_1_2___stage___block_6_clr;
_d___pip_5160_1_3___stage___block_6_clr = _q___pip_5160_1_3___stage___block_6_clr;
_d___pip_5160_1_4___stage___block_6_clr = _q___pip_5160_1_4___stage___block_6_clr;
_d___pip_5160_1_5___stage___block_6_clr = _q___pip_5160_1_5___stage___block_6_clr;
_d___pip_5160_1_6___stage___block_6_clr = _q___pip_5160_1_6___stage___block_6_clr;
_d___pip_5160_1_7___stage___block_6_clr = _q___pip_5160_1_7___stage___block_6_clr;
_d___pip_5160_1_8___stage___block_6_clr = _q___pip_5160_1_8___stage___block_6_clr;
_d___pip_5160_1_9___stage___block_6_clr = _q___pip_5160_1_9___stage___block_6_clr;
_d___pip_5160_1_10___stage___block_6_clr = _q___pip_5160_1_10___stage___block_6_clr;
_d___pip_5160_1_11___stage___block_6_clr = _q___pip_5160_1_11___stage___block_6_clr;
_d___pip_5160_1_12___stage___block_6_clr = _q___pip_5160_1_12___stage___block_6_clr;
_d___pip_5160_1_13___stage___block_6_clr = _q___pip_5160_1_13___stage___block_6_clr;
_d___pip_5160_1_14___stage___block_6_clr = _q___pip_5160_1_14___stage___block_6_clr;
_d___pip_5160_1_15___stage___block_6_clr = _q___pip_5160_1_15___stage___block_6_clr;
_d___pip_5160_1_16___stage___block_6_clr = _q___pip_5160_1_16___stage___block_6_clr;
_d___pip_5160_1_17___stage___block_6_clr = _q___pip_5160_1_17___stage___block_6_clr;
_d___pip_5160_1_18___stage___block_6_clr = _q___pip_5160_1_18___stage___block_6_clr;
_d___pip_5160_1_19___stage___block_6_clr = _q___pip_5160_1_19___stage___block_6_clr;
_d___pip_5160_1_20___stage___block_6_clr = _q___pip_5160_1_20___stage___block_6_clr;
_d___pip_5160_1_21___stage___block_6_clr = _q___pip_5160_1_21___stage___block_6_clr;
_d___pip_5160_1_22___stage___block_6_clr = _q___pip_5160_1_22___stage___block_6_clr;
_d___pip_5160_1_23___stage___block_6_clr = _q___pip_5160_1_23___stage___block_6_clr;
_d___pip_5160_1_24___stage___block_6_clr = _q___pip_5160_1_24___stage___block_6_clr;
_d___pip_5160_1_25___stage___block_6_clr = _q___pip_5160_1_25___stage___block_6_clr;
_d___pip_5160_1_26___stage___block_6_clr = _q___pip_5160_1_26___stage___block_6_clr;
_d___pip_5160_1_27___stage___block_6_clr = _q___pip_5160_1_27___stage___block_6_clr;
_d___pip_5160_1_28___stage___block_6_clr = _q___pip_5160_1_28___stage___block_6_clr;
_d___pip_5160_1_29___stage___block_6_clr = _q___pip_5160_1_29___stage___block_6_clr;
_d___pip_5160_1_30___stage___block_6_clr = _q___pip_5160_1_30___stage___block_6_clr;
_d___pip_5160_1_31___stage___block_6_clr = _q___pip_5160_1_31___stage___block_6_clr;
_d___pip_5160_1_32___stage___block_6_clr = _q___pip_5160_1_32___stage___block_6_clr;
_d___pip_5160_1_33___stage___block_6_clr = _q___pip_5160_1_33___stage___block_6_clr;
_d___pip_5160_1_34___stage___block_6_clr = _q___pip_5160_1_34___stage___block_6_clr;
_d___pip_5160_1_35___stage___block_6_clr = _q___pip_5160_1_35___stage___block_6_clr;
_d___pip_5160_1_36___stage___block_6_clr = _q___pip_5160_1_36___stage___block_6_clr;
_d___pip_5160_1_37___stage___block_6_clr = _q___pip_5160_1_37___stage___block_6_clr;
_d___pip_5160_1_38___stage___block_6_clr = _q___pip_5160_1_38___stage___block_6_clr;
_d___pip_5160_1_39___stage___block_6_clr = _q___pip_5160_1_39___stage___block_6_clr;
_d___pip_5160_1_40___stage___block_6_clr = _q___pip_5160_1_40___stage___block_6_clr;
_d___pip_5160_1_41___stage___block_6_clr = _q___pip_5160_1_41___stage___block_6_clr;
_d___pip_5160_1_42___stage___block_6_clr = _q___pip_5160_1_42___stage___block_6_clr;
_d___pip_5160_1_43___stage___block_6_clr = _q___pip_5160_1_43___stage___block_6_clr;
_d___pip_5160_1_44___stage___block_6_clr = _q___pip_5160_1_44___stage___block_6_clr;
_d___pip_5160_1_45___stage___block_6_clr = _q___pip_5160_1_45___stage___block_6_clr;
_d___pip_5160_1_46___stage___block_6_clr = _q___pip_5160_1_46___stage___block_6_clr;
_d___pip_5160_1_47___stage___block_6_clr = _q___pip_5160_1_47___stage___block_6_clr;
_d___pip_5160_1_48___stage___block_6_clr = _q___pip_5160_1_48___stage___block_6_clr;
_d___pip_5160_1_49___stage___block_6_clr = _q___pip_5160_1_49___stage___block_6_clr;
_d___pip_5160_1_50___stage___block_6_clr = _q___pip_5160_1_50___stage___block_6_clr;
_d___pip_5160_1_51___stage___block_6_clr = _q___pip_5160_1_51___stage___block_6_clr;
_d___pip_5160_1_52___stage___block_6_clr = _q___pip_5160_1_52___stage___block_6_clr;
_d___pip_5160_1_53___stage___block_6_clr = _q___pip_5160_1_53___stage___block_6_clr;
_d___pip_5160_1_54___stage___block_6_clr = _q___pip_5160_1_54___stage___block_6_clr;
_d___pip_5160_1_55___stage___block_6_clr = _q___pip_5160_1_55___stage___block_6_clr;
_d___pip_5160_1_56___stage___block_6_clr = _q___pip_5160_1_56___stage___block_6_clr;
_d___pip_5160_1_57___stage___block_6_clr = _q___pip_5160_1_57___stage___block_6_clr;
_d___pip_5160_1_58___stage___block_6_clr = _q___pip_5160_1_58___stage___block_6_clr;
_d___pip_5160_1_59___stage___block_6_clr = _q___pip_5160_1_59___stage___block_6_clr;
_d___pip_5160_1_60___stage___block_6_clr = _q___pip_5160_1_60___stage___block_6_clr;
_d___pip_5160_1_61___stage___block_6_clr = _q___pip_5160_1_61___stage___block_6_clr;
_d___pip_5160_1_62___stage___block_6_clr = _q___pip_5160_1_62___stage___block_6_clr;
_d___pip_5160_1_63___stage___block_6_clr = _q___pip_5160_1_63___stage___block_6_clr;
_d___pip_5160_1_64___stage___block_6_clr = _q___pip_5160_1_64___stage___block_6_clr;
_d___pip_5160_1_65___stage___block_6_clr = _q___pip_5160_1_65___stage___block_6_clr;
_d___pip_5160_1_66___stage___block_6_clr = _q___pip_5160_1_66___stage___block_6_clr;
_d___pip_5160_1_67___stage___block_6_clr = _q___pip_5160_1_67___stage___block_6_clr;
_d___pip_5160_1_68___stage___block_6_clr = _q___pip_5160_1_68___stage___block_6_clr;
_d___pip_5160_1_69___stage___block_6_clr = _q___pip_5160_1_69___stage___block_6_clr;
_d___pip_5160_1_70___stage___block_6_clr = _q___pip_5160_1_70___stage___block_6_clr;
_d___pip_5160_1_71___stage___block_6_clr = _q___pip_5160_1_71___stage___block_6_clr;
_d___pip_5160_1_72___stage___block_6_clr = _q___pip_5160_1_72___stage___block_6_clr;
_d___pip_5160_1_73___stage___block_6_clr = _q___pip_5160_1_73___stage___block_6_clr;
_d___pip_5160_1_74___stage___block_6_clr = _q___pip_5160_1_74___stage___block_6_clr;
_d___pip_5160_1_75___stage___block_6_clr = _q___pip_5160_1_75___stage___block_6_clr;
_d___pip_5160_1_76___stage___block_6_clr = _q___pip_5160_1_76___stage___block_6_clr;
_d___pip_5160_1_77___stage___block_6_clr = _q___pip_5160_1_77___stage___block_6_clr;
_d___pip_5160_1_78___stage___block_6_clr = _q___pip_5160_1_78___stage___block_6_clr;
_d___pip_5160_1_79___stage___block_6_clr = _q___pip_5160_1_79___stage___block_6_clr;
_d___pip_5160_1_80___stage___block_6_clr = _q___pip_5160_1_80___stage___block_6_clr;
_d___pip_5160_1_81___stage___block_6_clr = _q___pip_5160_1_81___stage___block_6_clr;
_d___pip_5160_1_82___stage___block_6_clr = _q___pip_5160_1_82___stage___block_6_clr;
_d___pip_5160_1_83___stage___block_6_clr = _q___pip_5160_1_83___stage___block_6_clr;
_d___pip_5160_1_84___stage___block_6_clr = _q___pip_5160_1_84___stage___block_6_clr;
_d___pip_5160_1_85___stage___block_6_clr = _q___pip_5160_1_85___stage___block_6_clr;
_d___pip_5160_1_86___stage___block_6_clr = _q___pip_5160_1_86___stage___block_6_clr;
_d___pip_5160_1_87___stage___block_6_clr = _q___pip_5160_1_87___stage___block_6_clr;
_d___pip_5160_1_88___stage___block_6_clr = _q___pip_5160_1_88___stage___block_6_clr;
_d___pip_5160_1_89___stage___block_6_clr = _q___pip_5160_1_89___stage___block_6_clr;
_d___pip_5160_1_90___stage___block_6_clr = _q___pip_5160_1_90___stage___block_6_clr;
_d___pip_5160_1_91___stage___block_6_clr = _q___pip_5160_1_91___stage___block_6_clr;
_d___pip_5160_1_92___stage___block_6_clr = _q___pip_5160_1_92___stage___block_6_clr;
_d___pip_5160_1_93___stage___block_6_clr = _q___pip_5160_1_93___stage___block_6_clr;
_d___pip_5160_1_94___stage___block_6_clr = _q___pip_5160_1_94___stage___block_6_clr;
_d___pip_5160_1_95___stage___block_6_clr = _q___pip_5160_1_95___stage___block_6_clr;
_d___pip_5160_1_96___stage___block_6_clr = _q___pip_5160_1_96___stage___block_6_clr;
_d___pip_5160_1_97___stage___block_6_clr = _q___pip_5160_1_97___stage___block_6_clr;
_d___pip_5160_1_98___stage___block_6_clr = _q___pip_5160_1_98___stage___block_6_clr;
_d___pip_5160_1_99___stage___block_6_clr = _q___pip_5160_1_99___stage___block_6_clr;
_d___pip_5160_1_100___stage___block_6_clr = _q___pip_5160_1_100___stage___block_6_clr;
_d___pip_5160_1_101___stage___block_6_clr = _q___pip_5160_1_101___stage___block_6_clr;
_d___pip_5160_1_102___stage___block_6_clr = _q___pip_5160_1_102___stage___block_6_clr;
_d___pip_5160_1_103___stage___block_6_clr = _q___pip_5160_1_103___stage___block_6_clr;
_d___pip_5160_1_104___stage___block_6_clr = _q___pip_5160_1_104___stage___block_6_clr;
_d___pip_5160_1_105___stage___block_6_clr = _q___pip_5160_1_105___stage___block_6_clr;
_d___pip_5160_1_106___stage___block_6_clr = _q___pip_5160_1_106___stage___block_6_clr;
_d___pip_5160_1_107___stage___block_6_clr = _q___pip_5160_1_107___stage___block_6_clr;
_d___pip_5160_1_108___stage___block_6_clr = _q___pip_5160_1_108___stage___block_6_clr;
_d___pip_5160_1_109___stage___block_6_clr = _q___pip_5160_1_109___stage___block_6_clr;
_d___pip_5160_1_110___stage___block_6_clr = _q___pip_5160_1_110___stage___block_6_clr;
_d___pip_5160_1_111___stage___block_6_clr = _q___pip_5160_1_111___stage___block_6_clr;
_d___pip_5160_1_112___stage___block_6_clr = _q___pip_5160_1_112___stage___block_6_clr;
_d___pip_5160_1_113___stage___block_6_clr = _q___pip_5160_1_113___stage___block_6_clr;
_d___pip_5160_1_114___stage___block_6_clr = _q___pip_5160_1_114___stage___block_6_clr;
_d___pip_5160_1_115___stage___block_6_clr = _q___pip_5160_1_115___stage___block_6_clr;
_d___pip_5160_1_116___stage___block_6_clr = _q___pip_5160_1_116___stage___block_6_clr;
_d___pip_5160_1_117___stage___block_6_clr = _q___pip_5160_1_117___stage___block_6_clr;
_d___pip_5160_1_118___stage___block_6_clr = _q___pip_5160_1_118___stage___block_6_clr;
_d___pip_5160_1_119___stage___block_6_clr = _q___pip_5160_1_119___stage___block_6_clr;
_d___pip_5160_1_120___stage___block_6_clr = _q___pip_5160_1_120___stage___block_6_clr;
_d___pip_5160_1_121___stage___block_6_clr = _q___pip_5160_1_121___stage___block_6_clr;
_d___pip_5160_1_122___stage___block_6_clr = _q___pip_5160_1_122___stage___block_6_clr;
_d___pip_5160_1_123___stage___block_6_clr = _q___pip_5160_1_123___stage___block_6_clr;
_d___pip_5160_1_124___stage___block_6_clr = _q___pip_5160_1_124___stage___block_6_clr;
_d___pip_5160_1_125___stage___block_6_clr = _q___pip_5160_1_125___stage___block_6_clr;
_d___pip_5160_1_126___stage___block_6_clr = _q___pip_5160_1_126___stage___block_6_clr;
_d___pip_5160_1_127___stage___block_6_clr = _q___pip_5160_1_127___stage___block_6_clr;
_d___pip_5160_1_128___stage___block_6_clr = _q___pip_5160_1_128___stage___block_6_clr;
_d___pip_5160_1_129___stage___block_6_clr = _q___pip_5160_1_129___stage___block_6_clr;
_d___pip_5160_1_130___stage___block_6_clr = _q___pip_5160_1_130___stage___block_6_clr;
_d___pip_5160_1_131___stage___block_6_clr = _q___pip_5160_1_131___stage___block_6_clr;
_d___pip_5160_1_132___stage___block_6_clr = _q___pip_5160_1_132___stage___block_6_clr;
_d___pip_5160_1_133___stage___block_6_clr = _q___pip_5160_1_133___stage___block_6_clr;
_d___pip_5160_1_134___stage___block_6_clr = _q___pip_5160_1_134___stage___block_6_clr;
_d___pip_5160_1_135___stage___block_6_clr = _q___pip_5160_1_135___stage___block_6_clr;
_d___pip_5160_1_0___stage___block_6_dist = _q___pip_5160_1_0___stage___block_6_dist;
_d___pip_5160_1_1___stage___block_6_dist = _q___pip_5160_1_1___stage___block_6_dist;
_d___pip_5160_1_2___stage___block_6_dist = _q___pip_5160_1_2___stage___block_6_dist;
_d___pip_5160_1_3___stage___block_6_dist = _q___pip_5160_1_3___stage___block_6_dist;
_d___pip_5160_1_4___stage___block_6_dist = _q___pip_5160_1_4___stage___block_6_dist;
_d___pip_5160_1_5___stage___block_6_dist = _q___pip_5160_1_5___stage___block_6_dist;
_d___pip_5160_1_6___stage___block_6_dist = _q___pip_5160_1_6___stage___block_6_dist;
_d___pip_5160_1_7___stage___block_6_dist = _q___pip_5160_1_7___stage___block_6_dist;
_d___pip_5160_1_8___stage___block_6_dist = _q___pip_5160_1_8___stage___block_6_dist;
_d___pip_5160_1_9___stage___block_6_dist = _q___pip_5160_1_9___stage___block_6_dist;
_d___pip_5160_1_10___stage___block_6_dist = _q___pip_5160_1_10___stage___block_6_dist;
_d___pip_5160_1_11___stage___block_6_dist = _q___pip_5160_1_11___stage___block_6_dist;
_d___pip_5160_1_12___stage___block_6_dist = _q___pip_5160_1_12___stage___block_6_dist;
_d___pip_5160_1_13___stage___block_6_dist = _q___pip_5160_1_13___stage___block_6_dist;
_d___pip_5160_1_14___stage___block_6_dist = _q___pip_5160_1_14___stage___block_6_dist;
_d___pip_5160_1_15___stage___block_6_dist = _q___pip_5160_1_15___stage___block_6_dist;
_d___pip_5160_1_16___stage___block_6_dist = _q___pip_5160_1_16___stage___block_6_dist;
_d___pip_5160_1_17___stage___block_6_dist = _q___pip_5160_1_17___stage___block_6_dist;
_d___pip_5160_1_18___stage___block_6_dist = _q___pip_5160_1_18___stage___block_6_dist;
_d___pip_5160_1_19___stage___block_6_dist = _q___pip_5160_1_19___stage___block_6_dist;
_d___pip_5160_1_20___stage___block_6_dist = _q___pip_5160_1_20___stage___block_6_dist;
_d___pip_5160_1_21___stage___block_6_dist = _q___pip_5160_1_21___stage___block_6_dist;
_d___pip_5160_1_22___stage___block_6_dist = _q___pip_5160_1_22___stage___block_6_dist;
_d___pip_5160_1_23___stage___block_6_dist = _q___pip_5160_1_23___stage___block_6_dist;
_d___pip_5160_1_24___stage___block_6_dist = _q___pip_5160_1_24___stage___block_6_dist;
_d___pip_5160_1_25___stage___block_6_dist = _q___pip_5160_1_25___stage___block_6_dist;
_d___pip_5160_1_26___stage___block_6_dist = _q___pip_5160_1_26___stage___block_6_dist;
_d___pip_5160_1_27___stage___block_6_dist = _q___pip_5160_1_27___stage___block_6_dist;
_d___pip_5160_1_28___stage___block_6_dist = _q___pip_5160_1_28___stage___block_6_dist;
_d___pip_5160_1_29___stage___block_6_dist = _q___pip_5160_1_29___stage___block_6_dist;
_d___pip_5160_1_30___stage___block_6_dist = _q___pip_5160_1_30___stage___block_6_dist;
_d___pip_5160_1_31___stage___block_6_dist = _q___pip_5160_1_31___stage___block_6_dist;
_d___pip_5160_1_32___stage___block_6_dist = _q___pip_5160_1_32___stage___block_6_dist;
_d___pip_5160_1_33___stage___block_6_dist = _q___pip_5160_1_33___stage___block_6_dist;
_d___pip_5160_1_34___stage___block_6_dist = _q___pip_5160_1_34___stage___block_6_dist;
_d___pip_5160_1_35___stage___block_6_dist = _q___pip_5160_1_35___stage___block_6_dist;
_d___pip_5160_1_36___stage___block_6_dist = _q___pip_5160_1_36___stage___block_6_dist;
_d___pip_5160_1_37___stage___block_6_dist = _q___pip_5160_1_37___stage___block_6_dist;
_d___pip_5160_1_38___stage___block_6_dist = _q___pip_5160_1_38___stage___block_6_dist;
_d___pip_5160_1_39___stage___block_6_dist = _q___pip_5160_1_39___stage___block_6_dist;
_d___pip_5160_1_40___stage___block_6_dist = _q___pip_5160_1_40___stage___block_6_dist;
_d___pip_5160_1_41___stage___block_6_dist = _q___pip_5160_1_41___stage___block_6_dist;
_d___pip_5160_1_42___stage___block_6_dist = _q___pip_5160_1_42___stage___block_6_dist;
_d___pip_5160_1_43___stage___block_6_dist = _q___pip_5160_1_43___stage___block_6_dist;
_d___pip_5160_1_44___stage___block_6_dist = _q___pip_5160_1_44___stage___block_6_dist;
_d___pip_5160_1_45___stage___block_6_dist = _q___pip_5160_1_45___stage___block_6_dist;
_d___pip_5160_1_46___stage___block_6_dist = _q___pip_5160_1_46___stage___block_6_dist;
_d___pip_5160_1_47___stage___block_6_dist = _q___pip_5160_1_47___stage___block_6_dist;
_d___pip_5160_1_48___stage___block_6_dist = _q___pip_5160_1_48___stage___block_6_dist;
_d___pip_5160_1_49___stage___block_6_dist = _q___pip_5160_1_49___stage___block_6_dist;
_d___pip_5160_1_50___stage___block_6_dist = _q___pip_5160_1_50___stage___block_6_dist;
_d___pip_5160_1_51___stage___block_6_dist = _q___pip_5160_1_51___stage___block_6_dist;
_d___pip_5160_1_52___stage___block_6_dist = _q___pip_5160_1_52___stage___block_6_dist;
_d___pip_5160_1_53___stage___block_6_dist = _q___pip_5160_1_53___stage___block_6_dist;
_d___pip_5160_1_54___stage___block_6_dist = _q___pip_5160_1_54___stage___block_6_dist;
_d___pip_5160_1_55___stage___block_6_dist = _q___pip_5160_1_55___stage___block_6_dist;
_d___pip_5160_1_56___stage___block_6_dist = _q___pip_5160_1_56___stage___block_6_dist;
_d___pip_5160_1_57___stage___block_6_dist = _q___pip_5160_1_57___stage___block_6_dist;
_d___pip_5160_1_58___stage___block_6_dist = _q___pip_5160_1_58___stage___block_6_dist;
_d___pip_5160_1_59___stage___block_6_dist = _q___pip_5160_1_59___stage___block_6_dist;
_d___pip_5160_1_60___stage___block_6_dist = _q___pip_5160_1_60___stage___block_6_dist;
_d___pip_5160_1_61___stage___block_6_dist = _q___pip_5160_1_61___stage___block_6_dist;
_d___pip_5160_1_62___stage___block_6_dist = _q___pip_5160_1_62___stage___block_6_dist;
_d___pip_5160_1_63___stage___block_6_dist = _q___pip_5160_1_63___stage___block_6_dist;
_d___pip_5160_1_64___stage___block_6_dist = _q___pip_5160_1_64___stage___block_6_dist;
_d___pip_5160_1_65___stage___block_6_dist = _q___pip_5160_1_65___stage___block_6_dist;
_d___pip_5160_1_66___stage___block_6_dist = _q___pip_5160_1_66___stage___block_6_dist;
_d___pip_5160_1_67___stage___block_6_dist = _q___pip_5160_1_67___stage___block_6_dist;
_d___pip_5160_1_68___stage___block_6_dist = _q___pip_5160_1_68___stage___block_6_dist;
_d___pip_5160_1_69___stage___block_6_dist = _q___pip_5160_1_69___stage___block_6_dist;
_d___pip_5160_1_70___stage___block_6_dist = _q___pip_5160_1_70___stage___block_6_dist;
_d___pip_5160_1_71___stage___block_6_dist = _q___pip_5160_1_71___stage___block_6_dist;
_d___pip_5160_1_72___stage___block_6_dist = _q___pip_5160_1_72___stage___block_6_dist;
_d___pip_5160_1_73___stage___block_6_dist = _q___pip_5160_1_73___stage___block_6_dist;
_d___pip_5160_1_74___stage___block_6_dist = _q___pip_5160_1_74___stage___block_6_dist;
_d___pip_5160_1_75___stage___block_6_dist = _q___pip_5160_1_75___stage___block_6_dist;
_d___pip_5160_1_76___stage___block_6_dist = _q___pip_5160_1_76___stage___block_6_dist;
_d___pip_5160_1_77___stage___block_6_dist = _q___pip_5160_1_77___stage___block_6_dist;
_d___pip_5160_1_78___stage___block_6_dist = _q___pip_5160_1_78___stage___block_6_dist;
_d___pip_5160_1_79___stage___block_6_dist = _q___pip_5160_1_79___stage___block_6_dist;
_d___pip_5160_1_80___stage___block_6_dist = _q___pip_5160_1_80___stage___block_6_dist;
_d___pip_5160_1_81___stage___block_6_dist = _q___pip_5160_1_81___stage___block_6_dist;
_d___pip_5160_1_82___stage___block_6_dist = _q___pip_5160_1_82___stage___block_6_dist;
_d___pip_5160_1_83___stage___block_6_dist = _q___pip_5160_1_83___stage___block_6_dist;
_d___pip_5160_1_84___stage___block_6_dist = _q___pip_5160_1_84___stage___block_6_dist;
_d___pip_5160_1_85___stage___block_6_dist = _q___pip_5160_1_85___stage___block_6_dist;
_d___pip_5160_1_86___stage___block_6_dist = _q___pip_5160_1_86___stage___block_6_dist;
_d___pip_5160_1_87___stage___block_6_dist = _q___pip_5160_1_87___stage___block_6_dist;
_d___pip_5160_1_88___stage___block_6_dist = _q___pip_5160_1_88___stage___block_6_dist;
_d___pip_5160_1_89___stage___block_6_dist = _q___pip_5160_1_89___stage___block_6_dist;
_d___pip_5160_1_90___stage___block_6_dist = _q___pip_5160_1_90___stage___block_6_dist;
_d___pip_5160_1_91___stage___block_6_dist = _q___pip_5160_1_91___stage___block_6_dist;
_d___pip_5160_1_92___stage___block_6_dist = _q___pip_5160_1_92___stage___block_6_dist;
_d___pip_5160_1_93___stage___block_6_dist = _q___pip_5160_1_93___stage___block_6_dist;
_d___pip_5160_1_94___stage___block_6_dist = _q___pip_5160_1_94___stage___block_6_dist;
_d___pip_5160_1_95___stage___block_6_dist = _q___pip_5160_1_95___stage___block_6_dist;
_d___pip_5160_1_96___stage___block_6_dist = _q___pip_5160_1_96___stage___block_6_dist;
_d___pip_5160_1_97___stage___block_6_dist = _q___pip_5160_1_97___stage___block_6_dist;
_d___pip_5160_1_98___stage___block_6_dist = _q___pip_5160_1_98___stage___block_6_dist;
_d___pip_5160_1_99___stage___block_6_dist = _q___pip_5160_1_99___stage___block_6_dist;
_d___pip_5160_1_100___stage___block_6_dist = _q___pip_5160_1_100___stage___block_6_dist;
_d___pip_5160_1_101___stage___block_6_dist = _q___pip_5160_1_101___stage___block_6_dist;
_d___pip_5160_1_102___stage___block_6_dist = _q___pip_5160_1_102___stage___block_6_dist;
_d___pip_5160_1_103___stage___block_6_dist = _q___pip_5160_1_103___stage___block_6_dist;
_d___pip_5160_1_104___stage___block_6_dist = _q___pip_5160_1_104___stage___block_6_dist;
_d___pip_5160_1_105___stage___block_6_dist = _q___pip_5160_1_105___stage___block_6_dist;
_d___pip_5160_1_106___stage___block_6_dist = _q___pip_5160_1_106___stage___block_6_dist;
_d___pip_5160_1_107___stage___block_6_dist = _q___pip_5160_1_107___stage___block_6_dist;
_d___pip_5160_1_108___stage___block_6_dist = _q___pip_5160_1_108___stage___block_6_dist;
_d___pip_5160_1_109___stage___block_6_dist = _q___pip_5160_1_109___stage___block_6_dist;
_d___pip_5160_1_110___stage___block_6_dist = _q___pip_5160_1_110___stage___block_6_dist;
_d___pip_5160_1_111___stage___block_6_dist = _q___pip_5160_1_111___stage___block_6_dist;
_d___pip_5160_1_112___stage___block_6_dist = _q___pip_5160_1_112___stage___block_6_dist;
_d___pip_5160_1_113___stage___block_6_dist = _q___pip_5160_1_113___stage___block_6_dist;
_d___pip_5160_1_114___stage___block_6_dist = _q___pip_5160_1_114___stage___block_6_dist;
_d___pip_5160_1_115___stage___block_6_dist = _q___pip_5160_1_115___stage___block_6_dist;
_d___pip_5160_1_116___stage___block_6_dist = _q___pip_5160_1_116___stage___block_6_dist;
_d___pip_5160_1_117___stage___block_6_dist = _q___pip_5160_1_117___stage___block_6_dist;
_d___pip_5160_1_118___stage___block_6_dist = _q___pip_5160_1_118___stage___block_6_dist;
_d___pip_5160_1_119___stage___block_6_dist = _q___pip_5160_1_119___stage___block_6_dist;
_d___pip_5160_1_120___stage___block_6_dist = _q___pip_5160_1_120___stage___block_6_dist;
_d___pip_5160_1_121___stage___block_6_dist = _q___pip_5160_1_121___stage___block_6_dist;
_d___pip_5160_1_122___stage___block_6_dist = _q___pip_5160_1_122___stage___block_6_dist;
_d___pip_5160_1_123___stage___block_6_dist = _q___pip_5160_1_123___stage___block_6_dist;
_d___pip_5160_1_124___stage___block_6_dist = _q___pip_5160_1_124___stage___block_6_dist;
_d___pip_5160_1_125___stage___block_6_dist = _q___pip_5160_1_125___stage___block_6_dist;
_d___pip_5160_1_126___stage___block_6_dist = _q___pip_5160_1_126___stage___block_6_dist;
_d___pip_5160_1_127___stage___block_6_dist = _q___pip_5160_1_127___stage___block_6_dist;
_d___pip_5160_1_128___stage___block_6_dist = _q___pip_5160_1_128___stage___block_6_dist;
_d___pip_5160_1_129___stage___block_6_dist = _q___pip_5160_1_129___stage___block_6_dist;
_d___pip_5160_1_130___stage___block_6_dist = _q___pip_5160_1_130___stage___block_6_dist;
_d___pip_5160_1_131___stage___block_6_dist = _q___pip_5160_1_131___stage___block_6_dist;
_d___pip_5160_1_132___stage___block_6_dist = _q___pip_5160_1_132___stage___block_6_dist;
_d___pip_5160_1_133___stage___block_6_dist = _q___pip_5160_1_133___stage___block_6_dist;
_d___pip_5160_1_134___stage___block_6_dist = _q___pip_5160_1_134___stage___block_6_dist;
_d___pip_5160_1_135___stage___block_6_dist = _q___pip_5160_1_135___stage___block_6_dist;
_d___pip_5160_1_0___stage___block_6_inside = _q___pip_5160_1_0___stage___block_6_inside;
_d___pip_5160_1_1___stage___block_6_inside = _q___pip_5160_1_1___stage___block_6_inside;
_d___pip_5160_1_2___stage___block_6_inside = _q___pip_5160_1_2___stage___block_6_inside;
_d___pip_5160_1_3___stage___block_6_inside = _q___pip_5160_1_3___stage___block_6_inside;
_d___pip_5160_1_4___stage___block_6_inside = _q___pip_5160_1_4___stage___block_6_inside;
_d___pip_5160_1_5___stage___block_6_inside = _q___pip_5160_1_5___stage___block_6_inside;
_d___pip_5160_1_6___stage___block_6_inside = _q___pip_5160_1_6___stage___block_6_inside;
_d___pip_5160_1_7___stage___block_6_inside = _q___pip_5160_1_7___stage___block_6_inside;
_d___pip_5160_1_8___stage___block_6_inside = _q___pip_5160_1_8___stage___block_6_inside;
_d___pip_5160_1_9___stage___block_6_inside = _q___pip_5160_1_9___stage___block_6_inside;
_d___pip_5160_1_10___stage___block_6_inside = _q___pip_5160_1_10___stage___block_6_inside;
_d___pip_5160_1_11___stage___block_6_inside = _q___pip_5160_1_11___stage___block_6_inside;
_d___pip_5160_1_12___stage___block_6_inside = _q___pip_5160_1_12___stage___block_6_inside;
_d___pip_5160_1_13___stage___block_6_inside = _q___pip_5160_1_13___stage___block_6_inside;
_d___pip_5160_1_14___stage___block_6_inside = _q___pip_5160_1_14___stage___block_6_inside;
_d___pip_5160_1_15___stage___block_6_inside = _q___pip_5160_1_15___stage___block_6_inside;
_d___pip_5160_1_16___stage___block_6_inside = _q___pip_5160_1_16___stage___block_6_inside;
_d___pip_5160_1_17___stage___block_6_inside = _q___pip_5160_1_17___stage___block_6_inside;
_d___pip_5160_1_18___stage___block_6_inside = _q___pip_5160_1_18___stage___block_6_inside;
_d___pip_5160_1_19___stage___block_6_inside = _q___pip_5160_1_19___stage___block_6_inside;
_d___pip_5160_1_20___stage___block_6_inside = _q___pip_5160_1_20___stage___block_6_inside;
_d___pip_5160_1_21___stage___block_6_inside = _q___pip_5160_1_21___stage___block_6_inside;
_d___pip_5160_1_22___stage___block_6_inside = _q___pip_5160_1_22___stage___block_6_inside;
_d___pip_5160_1_23___stage___block_6_inside = _q___pip_5160_1_23___stage___block_6_inside;
_d___pip_5160_1_24___stage___block_6_inside = _q___pip_5160_1_24___stage___block_6_inside;
_d___pip_5160_1_25___stage___block_6_inside = _q___pip_5160_1_25___stage___block_6_inside;
_d___pip_5160_1_26___stage___block_6_inside = _q___pip_5160_1_26___stage___block_6_inside;
_d___pip_5160_1_27___stage___block_6_inside = _q___pip_5160_1_27___stage___block_6_inside;
_d___pip_5160_1_28___stage___block_6_inside = _q___pip_5160_1_28___stage___block_6_inside;
_d___pip_5160_1_29___stage___block_6_inside = _q___pip_5160_1_29___stage___block_6_inside;
_d___pip_5160_1_30___stage___block_6_inside = _q___pip_5160_1_30___stage___block_6_inside;
_d___pip_5160_1_31___stage___block_6_inside = _q___pip_5160_1_31___stage___block_6_inside;
_d___pip_5160_1_32___stage___block_6_inside = _q___pip_5160_1_32___stage___block_6_inside;
_d___pip_5160_1_33___stage___block_6_inside = _q___pip_5160_1_33___stage___block_6_inside;
_d___pip_5160_1_34___stage___block_6_inside = _q___pip_5160_1_34___stage___block_6_inside;
_d___pip_5160_1_35___stage___block_6_inside = _q___pip_5160_1_35___stage___block_6_inside;
_d___pip_5160_1_36___stage___block_6_inside = _q___pip_5160_1_36___stage___block_6_inside;
_d___pip_5160_1_37___stage___block_6_inside = _q___pip_5160_1_37___stage___block_6_inside;
_d___pip_5160_1_38___stage___block_6_inside = _q___pip_5160_1_38___stage___block_6_inside;
_d___pip_5160_1_39___stage___block_6_inside = _q___pip_5160_1_39___stage___block_6_inside;
_d___pip_5160_1_40___stage___block_6_inside = _q___pip_5160_1_40___stage___block_6_inside;
_d___pip_5160_1_41___stage___block_6_inside = _q___pip_5160_1_41___stage___block_6_inside;
_d___pip_5160_1_42___stage___block_6_inside = _q___pip_5160_1_42___stage___block_6_inside;
_d___pip_5160_1_43___stage___block_6_inside = _q___pip_5160_1_43___stage___block_6_inside;
_d___pip_5160_1_44___stage___block_6_inside = _q___pip_5160_1_44___stage___block_6_inside;
_d___pip_5160_1_45___stage___block_6_inside = _q___pip_5160_1_45___stage___block_6_inside;
_d___pip_5160_1_46___stage___block_6_inside = _q___pip_5160_1_46___stage___block_6_inside;
_d___pip_5160_1_47___stage___block_6_inside = _q___pip_5160_1_47___stage___block_6_inside;
_d___pip_5160_1_48___stage___block_6_inside = _q___pip_5160_1_48___stage___block_6_inside;
_d___pip_5160_1_49___stage___block_6_inside = _q___pip_5160_1_49___stage___block_6_inside;
_d___pip_5160_1_50___stage___block_6_inside = _q___pip_5160_1_50___stage___block_6_inside;
_d___pip_5160_1_51___stage___block_6_inside = _q___pip_5160_1_51___stage___block_6_inside;
_d___pip_5160_1_52___stage___block_6_inside = _q___pip_5160_1_52___stage___block_6_inside;
_d___pip_5160_1_53___stage___block_6_inside = _q___pip_5160_1_53___stage___block_6_inside;
_d___pip_5160_1_54___stage___block_6_inside = _q___pip_5160_1_54___stage___block_6_inside;
_d___pip_5160_1_55___stage___block_6_inside = _q___pip_5160_1_55___stage___block_6_inside;
_d___pip_5160_1_56___stage___block_6_inside = _q___pip_5160_1_56___stage___block_6_inside;
_d___pip_5160_1_57___stage___block_6_inside = _q___pip_5160_1_57___stage___block_6_inside;
_d___pip_5160_1_58___stage___block_6_inside = _q___pip_5160_1_58___stage___block_6_inside;
_d___pip_5160_1_59___stage___block_6_inside = _q___pip_5160_1_59___stage___block_6_inside;
_d___pip_5160_1_60___stage___block_6_inside = _q___pip_5160_1_60___stage___block_6_inside;
_d___pip_5160_1_61___stage___block_6_inside = _q___pip_5160_1_61___stage___block_6_inside;
_d___pip_5160_1_62___stage___block_6_inside = _q___pip_5160_1_62___stage___block_6_inside;
_d___pip_5160_1_63___stage___block_6_inside = _q___pip_5160_1_63___stage___block_6_inside;
_d___pip_5160_1_64___stage___block_6_inside = _q___pip_5160_1_64___stage___block_6_inside;
_d___pip_5160_1_65___stage___block_6_inside = _q___pip_5160_1_65___stage___block_6_inside;
_d___pip_5160_1_66___stage___block_6_inside = _q___pip_5160_1_66___stage___block_6_inside;
_d___pip_5160_1_67___stage___block_6_inside = _q___pip_5160_1_67___stage___block_6_inside;
_d___pip_5160_1_68___stage___block_6_inside = _q___pip_5160_1_68___stage___block_6_inside;
_d___pip_5160_1_69___stage___block_6_inside = _q___pip_5160_1_69___stage___block_6_inside;
_d___pip_5160_1_70___stage___block_6_inside = _q___pip_5160_1_70___stage___block_6_inside;
_d___pip_5160_1_71___stage___block_6_inside = _q___pip_5160_1_71___stage___block_6_inside;
_d___pip_5160_1_72___stage___block_6_inside = _q___pip_5160_1_72___stage___block_6_inside;
_d___pip_5160_1_73___stage___block_6_inside = _q___pip_5160_1_73___stage___block_6_inside;
_d___pip_5160_1_74___stage___block_6_inside = _q___pip_5160_1_74___stage___block_6_inside;
_d___pip_5160_1_75___stage___block_6_inside = _q___pip_5160_1_75___stage___block_6_inside;
_d___pip_5160_1_76___stage___block_6_inside = _q___pip_5160_1_76___stage___block_6_inside;
_d___pip_5160_1_77___stage___block_6_inside = _q___pip_5160_1_77___stage___block_6_inside;
_d___pip_5160_1_78___stage___block_6_inside = _q___pip_5160_1_78___stage___block_6_inside;
_d___pip_5160_1_79___stage___block_6_inside = _q___pip_5160_1_79___stage___block_6_inside;
_d___pip_5160_1_80___stage___block_6_inside = _q___pip_5160_1_80___stage___block_6_inside;
_d___pip_5160_1_81___stage___block_6_inside = _q___pip_5160_1_81___stage___block_6_inside;
_d___pip_5160_1_82___stage___block_6_inside = _q___pip_5160_1_82___stage___block_6_inside;
_d___pip_5160_1_83___stage___block_6_inside = _q___pip_5160_1_83___stage___block_6_inside;
_d___pip_5160_1_84___stage___block_6_inside = _q___pip_5160_1_84___stage___block_6_inside;
_d___pip_5160_1_85___stage___block_6_inside = _q___pip_5160_1_85___stage___block_6_inside;
_d___pip_5160_1_86___stage___block_6_inside = _q___pip_5160_1_86___stage___block_6_inside;
_d___pip_5160_1_87___stage___block_6_inside = _q___pip_5160_1_87___stage___block_6_inside;
_d___pip_5160_1_88___stage___block_6_inside = _q___pip_5160_1_88___stage___block_6_inside;
_d___pip_5160_1_89___stage___block_6_inside = _q___pip_5160_1_89___stage___block_6_inside;
_d___pip_5160_1_90___stage___block_6_inside = _q___pip_5160_1_90___stage___block_6_inside;
_d___pip_5160_1_91___stage___block_6_inside = _q___pip_5160_1_91___stage___block_6_inside;
_d___pip_5160_1_92___stage___block_6_inside = _q___pip_5160_1_92___stage___block_6_inside;
_d___pip_5160_1_93___stage___block_6_inside = _q___pip_5160_1_93___stage___block_6_inside;
_d___pip_5160_1_94___stage___block_6_inside = _q___pip_5160_1_94___stage___block_6_inside;
_d___pip_5160_1_95___stage___block_6_inside = _q___pip_5160_1_95___stage___block_6_inside;
_d___pip_5160_1_96___stage___block_6_inside = _q___pip_5160_1_96___stage___block_6_inside;
_d___pip_5160_1_97___stage___block_6_inside = _q___pip_5160_1_97___stage___block_6_inside;
_d___pip_5160_1_98___stage___block_6_inside = _q___pip_5160_1_98___stage___block_6_inside;
_d___pip_5160_1_99___stage___block_6_inside = _q___pip_5160_1_99___stage___block_6_inside;
_d___pip_5160_1_100___stage___block_6_inside = _q___pip_5160_1_100___stage___block_6_inside;
_d___pip_5160_1_101___stage___block_6_inside = _q___pip_5160_1_101___stage___block_6_inside;
_d___pip_5160_1_102___stage___block_6_inside = _q___pip_5160_1_102___stage___block_6_inside;
_d___pip_5160_1_103___stage___block_6_inside = _q___pip_5160_1_103___stage___block_6_inside;
_d___pip_5160_1_104___stage___block_6_inside = _q___pip_5160_1_104___stage___block_6_inside;
_d___pip_5160_1_105___stage___block_6_inside = _q___pip_5160_1_105___stage___block_6_inside;
_d___pip_5160_1_106___stage___block_6_inside = _q___pip_5160_1_106___stage___block_6_inside;
_d___pip_5160_1_107___stage___block_6_inside = _q___pip_5160_1_107___stage___block_6_inside;
_d___pip_5160_1_108___stage___block_6_inside = _q___pip_5160_1_108___stage___block_6_inside;
_d___pip_5160_1_109___stage___block_6_inside = _q___pip_5160_1_109___stage___block_6_inside;
_d___pip_5160_1_110___stage___block_6_inside = _q___pip_5160_1_110___stage___block_6_inside;
_d___pip_5160_1_111___stage___block_6_inside = _q___pip_5160_1_111___stage___block_6_inside;
_d___pip_5160_1_112___stage___block_6_inside = _q___pip_5160_1_112___stage___block_6_inside;
_d___pip_5160_1_113___stage___block_6_inside = _q___pip_5160_1_113___stage___block_6_inside;
_d___pip_5160_1_114___stage___block_6_inside = _q___pip_5160_1_114___stage___block_6_inside;
_d___pip_5160_1_115___stage___block_6_inside = _q___pip_5160_1_115___stage___block_6_inside;
_d___pip_5160_1_116___stage___block_6_inside = _q___pip_5160_1_116___stage___block_6_inside;
_d___pip_5160_1_117___stage___block_6_inside = _q___pip_5160_1_117___stage___block_6_inside;
_d___pip_5160_1_118___stage___block_6_inside = _q___pip_5160_1_118___stage___block_6_inside;
_d___pip_5160_1_119___stage___block_6_inside = _q___pip_5160_1_119___stage___block_6_inside;
_d___pip_5160_1_120___stage___block_6_inside = _q___pip_5160_1_120___stage___block_6_inside;
_d___pip_5160_1_121___stage___block_6_inside = _q___pip_5160_1_121___stage___block_6_inside;
_d___pip_5160_1_122___stage___block_6_inside = _q___pip_5160_1_122___stage___block_6_inside;
_d___pip_5160_1_123___stage___block_6_inside = _q___pip_5160_1_123___stage___block_6_inside;
_d___pip_5160_1_124___stage___block_6_inside = _q___pip_5160_1_124___stage___block_6_inside;
_d___pip_5160_1_125___stage___block_6_inside = _q___pip_5160_1_125___stage___block_6_inside;
_d___pip_5160_1_126___stage___block_6_inside = _q___pip_5160_1_126___stage___block_6_inside;
_d___pip_5160_1_127___stage___block_6_inside = _q___pip_5160_1_127___stage___block_6_inside;
_d___pip_5160_1_128___stage___block_6_inside = _q___pip_5160_1_128___stage___block_6_inside;
_d___pip_5160_1_129___stage___block_6_inside = _q___pip_5160_1_129___stage___block_6_inside;
_d___pip_5160_1_130___stage___block_6_inside = _q___pip_5160_1_130___stage___block_6_inside;
_d___pip_5160_1_131___stage___block_6_inside = _q___pip_5160_1_131___stage___block_6_inside;
_d___pip_5160_1_132___stage___block_6_inside = _q___pip_5160_1_132___stage___block_6_inside;
_d___pip_5160_1_133___stage___block_6_inside = _q___pip_5160_1_133___stage___block_6_inside;
_d___pip_5160_1_134___stage___block_6_inside = _q___pip_5160_1_134___stage___block_6_inside;
_d___pip_5160_1_0___stage___block_6_view_x = _q___pip_5160_1_0___stage___block_6_view_x;
_d___pip_5160_1_1___stage___block_6_view_x = _q___pip_5160_1_1___stage___block_6_view_x;
_d___pip_5160_1_2___stage___block_6_view_x = _q___pip_5160_1_2___stage___block_6_view_x;
_d___pip_5160_1_3___stage___block_6_view_x = _q___pip_5160_1_3___stage___block_6_view_x;
_d___pip_5160_1_0___stage___block_6_view_y = _q___pip_5160_1_0___stage___block_6_view_y;
_d___pip_5160_1_1___stage___block_6_view_y = _q___pip_5160_1_1___stage___block_6_view_y;
_d___pip_5160_1_2___stage___block_6_view_y = _q___pip_5160_1_2___stage___block_6_view_y;
_d___pip_5160_1_3___stage___block_6_view_y = _q___pip_5160_1_3___stage___block_6_view_y;
_d___pip_5160_1_4___stage___block_6_view_y = _q___pip_5160_1_4___stage___block_6_view_y;
_d___pip_5160_1_0___stage___block_6_view_z = _q___pip_5160_1_0___stage___block_6_view_z;
_d___pip_5160_1_1___stage___block_6_view_z = _q___pip_5160_1_1___stage___block_6_view_z;
_d___pip_5160_1_2___stage___block_6_view_z = _q___pip_5160_1_2___stage___block_6_view_z;
_d___pip_5160_1_3___stage___block_6_view_z = _q___pip_5160_1_3___stage___block_6_view_z;
_d___pip_5160_1_0___stage___block_6_vxsz = _q___pip_5160_1_0___stage___block_6_vxsz;
_d___pip_5160_1_1___stage___block_6_vxsz = _q___pip_5160_1_1___stage___block_6_vxsz;
_d___pip_5160_1_2___stage___block_6_vxsz = _q___pip_5160_1_2___stage___block_6_vxsz;
_d___pip_5160_1_3___stage___block_6_vxsz = _q___pip_5160_1_3___stage___block_6_vxsz;
_d___pip_5160_1_4___stage___block_6_vxsz = _q___pip_5160_1_4___stage___block_6_vxsz;
_d___pip_5160_1_5___stage___block_6_vxsz = _q___pip_5160_1_5___stage___block_6_vxsz;
_d___pip_5160_1_6___stage___block_6_vxsz = _q___pip_5160_1_6___stage___block_6_vxsz;
_d___pip_5160_1_1___stage___block_7_cs0 = _q___pip_5160_1_1___stage___block_7_cs0;
_d___pip_5160_1_2___stage___block_7_cs0 = _q___pip_5160_1_2___stage___block_7_cs0;
_d___pip_5160_1_3___stage___block_7_cs0 = _q___pip_5160_1_3___stage___block_7_cs0;
_d___pip_5160_1_1___stage___block_7_ss0 = _q___pip_5160_1_1___stage___block_7_ss0;
_d___pip_5160_1_2___stage___block_7_ss0 = _q___pip_5160_1_2___stage___block_7_ss0;
_d___pip_5160_1_3___stage___block_7_ss0 = _q___pip_5160_1_3___stage___block_7_ss0;
_d_pix_r = _q_pix_r;
_d_pix_g = _q_pix_g;
_d_pix_b = _q_pix_b;
_d__idx_fsm0 = _q__idx_fsm0;
_d__idx_fsm___pip_5160_1_0 = _q__idx_fsm___pip_5160_1_0;
_d__full_fsm___pip_5160_1_0 = _q__full_fsm___pip_5160_1_0;
_t__stall_fsm___pip_5160_1_0 = 0;
_t__1stdisable_fsm___pip_5160_1_0 = 0;
_d__idx_fsm___pip_5160_1_1 = _q__idx_fsm___pip_5160_1_1;
_d__full_fsm___pip_5160_1_1 = _q__full_fsm___pip_5160_1_1;
_t__stall_fsm___pip_5160_1_1 = 0;
_t__1stdisable_fsm___pip_5160_1_1 = 0;
_d__idx_fsm___pip_5160_1_2 = _q__idx_fsm___pip_5160_1_2;
_d__full_fsm___pip_5160_1_2 = _q__full_fsm___pip_5160_1_2;
_t__stall_fsm___pip_5160_1_2 = 0;
_t__1stdisable_fsm___pip_5160_1_2 = 0;
_d__idx_fsm___pip_5160_1_3 = _q__idx_fsm___pip_5160_1_3;
_d__full_fsm___pip_5160_1_3 = _q__full_fsm___pip_5160_1_3;
_t__stall_fsm___pip_5160_1_3 = 0;
_t__1stdisable_fsm___pip_5160_1_3 = 0;
_d__idx_fsm___pip_5160_1_4 = _q__idx_fsm___pip_5160_1_4;
_d__full_fsm___pip_5160_1_4 = _q__full_fsm___pip_5160_1_4;
_t__stall_fsm___pip_5160_1_4 = 0;
_t__1stdisable_fsm___pip_5160_1_4 = 0;
_d__idx_fsm___pip_5160_1_5 = _q__idx_fsm___pip_5160_1_5;
_d__full_fsm___pip_5160_1_5 = _q__full_fsm___pip_5160_1_5;
_t__stall_fsm___pip_5160_1_5 = 0;
_t__1stdisable_fsm___pip_5160_1_5 = 0;
_d__idx_fsm___pip_5160_1_6 = _q__idx_fsm___pip_5160_1_6;
_d__full_fsm___pip_5160_1_6 = _q__full_fsm___pip_5160_1_6;
_t__stall_fsm___pip_5160_1_6 = 0;
_t__1stdisable_fsm___pip_5160_1_6 = 0;
_d__idx_fsm___pip_5160_1_7 = _q__idx_fsm___pip_5160_1_7;
_d__full_fsm___pip_5160_1_7 = _q__full_fsm___pip_5160_1_7;
_t__stall_fsm___pip_5160_1_7 = 0;
_t__1stdisable_fsm___pip_5160_1_7 = 0;
_d__idx_fsm___pip_5160_1_8 = _q__idx_fsm___pip_5160_1_8;
_d__full_fsm___pip_5160_1_8 = _q__full_fsm___pip_5160_1_8;
_t__stall_fsm___pip_5160_1_8 = 0;
_t__1stdisable_fsm___pip_5160_1_8 = 0;
_d__idx_fsm___pip_5160_1_9 = _q__idx_fsm___pip_5160_1_9;
_d__full_fsm___pip_5160_1_9 = _q__full_fsm___pip_5160_1_9;
_t__stall_fsm___pip_5160_1_9 = 0;
_t__1stdisable_fsm___pip_5160_1_9 = 0;
_d__idx_fsm___pip_5160_1_10 = _q__idx_fsm___pip_5160_1_10;
_d__full_fsm___pip_5160_1_10 = _q__full_fsm___pip_5160_1_10;
_t__stall_fsm___pip_5160_1_10 = 0;
_t__1stdisable_fsm___pip_5160_1_10 = 0;
_d__idx_fsm___pip_5160_1_11 = _q__idx_fsm___pip_5160_1_11;
_d__full_fsm___pip_5160_1_11 = _q__full_fsm___pip_5160_1_11;
_t__stall_fsm___pip_5160_1_11 = 0;
_t__1stdisable_fsm___pip_5160_1_11 = 0;
_d__idx_fsm___pip_5160_1_12 = _q__idx_fsm___pip_5160_1_12;
_d__full_fsm___pip_5160_1_12 = _q__full_fsm___pip_5160_1_12;
_t__stall_fsm___pip_5160_1_12 = 0;
_t__1stdisable_fsm___pip_5160_1_12 = 0;
_d__idx_fsm___pip_5160_1_13 = _q__idx_fsm___pip_5160_1_13;
_d__full_fsm___pip_5160_1_13 = _q__full_fsm___pip_5160_1_13;
_t__stall_fsm___pip_5160_1_13 = 0;
_t__1stdisable_fsm___pip_5160_1_13 = 0;
_d__idx_fsm___pip_5160_1_14 = _q__idx_fsm___pip_5160_1_14;
_d__full_fsm___pip_5160_1_14 = _q__full_fsm___pip_5160_1_14;
_t__stall_fsm___pip_5160_1_14 = 0;
_t__1stdisable_fsm___pip_5160_1_14 = 0;
_d__idx_fsm___pip_5160_1_15 = _q__idx_fsm___pip_5160_1_15;
_d__full_fsm___pip_5160_1_15 = _q__full_fsm___pip_5160_1_15;
_t__stall_fsm___pip_5160_1_15 = 0;
_t__1stdisable_fsm___pip_5160_1_15 = 0;
_d__idx_fsm___pip_5160_1_16 = _q__idx_fsm___pip_5160_1_16;
_d__full_fsm___pip_5160_1_16 = _q__full_fsm___pip_5160_1_16;
_t__stall_fsm___pip_5160_1_16 = 0;
_t__1stdisable_fsm___pip_5160_1_16 = 0;
_d__idx_fsm___pip_5160_1_17 = _q__idx_fsm___pip_5160_1_17;
_d__full_fsm___pip_5160_1_17 = _q__full_fsm___pip_5160_1_17;
_t__stall_fsm___pip_5160_1_17 = 0;
_t__1stdisable_fsm___pip_5160_1_17 = 0;
_d__idx_fsm___pip_5160_1_18 = _q__idx_fsm___pip_5160_1_18;
_d__full_fsm___pip_5160_1_18 = _q__full_fsm___pip_5160_1_18;
_t__stall_fsm___pip_5160_1_18 = 0;
_t__1stdisable_fsm___pip_5160_1_18 = 0;
_d__idx_fsm___pip_5160_1_19 = _q__idx_fsm___pip_5160_1_19;
_d__full_fsm___pip_5160_1_19 = _q__full_fsm___pip_5160_1_19;
_t__stall_fsm___pip_5160_1_19 = 0;
_t__1stdisable_fsm___pip_5160_1_19 = 0;
_d__idx_fsm___pip_5160_1_20 = _q__idx_fsm___pip_5160_1_20;
_d__full_fsm___pip_5160_1_20 = _q__full_fsm___pip_5160_1_20;
_t__stall_fsm___pip_5160_1_20 = 0;
_t__1stdisable_fsm___pip_5160_1_20 = 0;
_d__idx_fsm___pip_5160_1_21 = _q__idx_fsm___pip_5160_1_21;
_d__full_fsm___pip_5160_1_21 = _q__full_fsm___pip_5160_1_21;
_t__stall_fsm___pip_5160_1_21 = 0;
_t__1stdisable_fsm___pip_5160_1_21 = 0;
_d__idx_fsm___pip_5160_1_22 = _q__idx_fsm___pip_5160_1_22;
_d__full_fsm___pip_5160_1_22 = _q__full_fsm___pip_5160_1_22;
_t__stall_fsm___pip_5160_1_22 = 0;
_t__1stdisable_fsm___pip_5160_1_22 = 0;
_d__idx_fsm___pip_5160_1_23 = _q__idx_fsm___pip_5160_1_23;
_d__full_fsm___pip_5160_1_23 = _q__full_fsm___pip_5160_1_23;
_t__stall_fsm___pip_5160_1_23 = 0;
_t__1stdisable_fsm___pip_5160_1_23 = 0;
_d__idx_fsm___pip_5160_1_24 = _q__idx_fsm___pip_5160_1_24;
_d__full_fsm___pip_5160_1_24 = _q__full_fsm___pip_5160_1_24;
_t__stall_fsm___pip_5160_1_24 = 0;
_t__1stdisable_fsm___pip_5160_1_24 = 0;
_d__idx_fsm___pip_5160_1_25 = _q__idx_fsm___pip_5160_1_25;
_d__full_fsm___pip_5160_1_25 = _q__full_fsm___pip_5160_1_25;
_t__stall_fsm___pip_5160_1_25 = 0;
_t__1stdisable_fsm___pip_5160_1_25 = 0;
_d__idx_fsm___pip_5160_1_26 = _q__idx_fsm___pip_5160_1_26;
_d__full_fsm___pip_5160_1_26 = _q__full_fsm___pip_5160_1_26;
_t__stall_fsm___pip_5160_1_26 = 0;
_t__1stdisable_fsm___pip_5160_1_26 = 0;
_d__idx_fsm___pip_5160_1_27 = _q__idx_fsm___pip_5160_1_27;
_d__full_fsm___pip_5160_1_27 = _q__full_fsm___pip_5160_1_27;
_t__stall_fsm___pip_5160_1_27 = 0;
_t__1stdisable_fsm___pip_5160_1_27 = 0;
_d__idx_fsm___pip_5160_1_28 = _q__idx_fsm___pip_5160_1_28;
_d__full_fsm___pip_5160_1_28 = _q__full_fsm___pip_5160_1_28;
_t__stall_fsm___pip_5160_1_28 = 0;
_t__1stdisable_fsm___pip_5160_1_28 = 0;
_d__idx_fsm___pip_5160_1_29 = _q__idx_fsm___pip_5160_1_29;
_d__full_fsm___pip_5160_1_29 = _q__full_fsm___pip_5160_1_29;
_t__stall_fsm___pip_5160_1_29 = 0;
_t__1stdisable_fsm___pip_5160_1_29 = 0;
_d__idx_fsm___pip_5160_1_30 = _q__idx_fsm___pip_5160_1_30;
_d__full_fsm___pip_5160_1_30 = _q__full_fsm___pip_5160_1_30;
_t__stall_fsm___pip_5160_1_30 = 0;
_t__1stdisable_fsm___pip_5160_1_30 = 0;
_d__idx_fsm___pip_5160_1_31 = _q__idx_fsm___pip_5160_1_31;
_d__full_fsm___pip_5160_1_31 = _q__full_fsm___pip_5160_1_31;
_t__stall_fsm___pip_5160_1_31 = 0;
_t__1stdisable_fsm___pip_5160_1_31 = 0;
_d__idx_fsm___pip_5160_1_32 = _q__idx_fsm___pip_5160_1_32;
_d__full_fsm___pip_5160_1_32 = _q__full_fsm___pip_5160_1_32;
_t__stall_fsm___pip_5160_1_32 = 0;
_t__1stdisable_fsm___pip_5160_1_32 = 0;
_d__idx_fsm___pip_5160_1_33 = _q__idx_fsm___pip_5160_1_33;
_d__full_fsm___pip_5160_1_33 = _q__full_fsm___pip_5160_1_33;
_t__stall_fsm___pip_5160_1_33 = 0;
_t__1stdisable_fsm___pip_5160_1_33 = 0;
_d__idx_fsm___pip_5160_1_34 = _q__idx_fsm___pip_5160_1_34;
_d__full_fsm___pip_5160_1_34 = _q__full_fsm___pip_5160_1_34;
_t__stall_fsm___pip_5160_1_34 = 0;
_t__1stdisable_fsm___pip_5160_1_34 = 0;
_d__idx_fsm___pip_5160_1_35 = _q__idx_fsm___pip_5160_1_35;
_d__full_fsm___pip_5160_1_35 = _q__full_fsm___pip_5160_1_35;
_t__stall_fsm___pip_5160_1_35 = 0;
_t__1stdisable_fsm___pip_5160_1_35 = 0;
_d__idx_fsm___pip_5160_1_36 = _q__idx_fsm___pip_5160_1_36;
_d__full_fsm___pip_5160_1_36 = _q__full_fsm___pip_5160_1_36;
_t__stall_fsm___pip_5160_1_36 = 0;
_t__1stdisable_fsm___pip_5160_1_36 = 0;
_d__idx_fsm___pip_5160_1_37 = _q__idx_fsm___pip_5160_1_37;
_d__full_fsm___pip_5160_1_37 = _q__full_fsm___pip_5160_1_37;
_t__stall_fsm___pip_5160_1_37 = 0;
_t__1stdisable_fsm___pip_5160_1_37 = 0;
_d__idx_fsm___pip_5160_1_38 = _q__idx_fsm___pip_5160_1_38;
_d__full_fsm___pip_5160_1_38 = _q__full_fsm___pip_5160_1_38;
_t__stall_fsm___pip_5160_1_38 = 0;
_t__1stdisable_fsm___pip_5160_1_38 = 0;
_d__idx_fsm___pip_5160_1_39 = _q__idx_fsm___pip_5160_1_39;
_d__full_fsm___pip_5160_1_39 = _q__full_fsm___pip_5160_1_39;
_t__stall_fsm___pip_5160_1_39 = 0;
_t__1stdisable_fsm___pip_5160_1_39 = 0;
_d__idx_fsm___pip_5160_1_40 = _q__idx_fsm___pip_5160_1_40;
_d__full_fsm___pip_5160_1_40 = _q__full_fsm___pip_5160_1_40;
_t__stall_fsm___pip_5160_1_40 = 0;
_t__1stdisable_fsm___pip_5160_1_40 = 0;
_d__idx_fsm___pip_5160_1_41 = _q__idx_fsm___pip_5160_1_41;
_d__full_fsm___pip_5160_1_41 = _q__full_fsm___pip_5160_1_41;
_t__stall_fsm___pip_5160_1_41 = 0;
_t__1stdisable_fsm___pip_5160_1_41 = 0;
_d__idx_fsm___pip_5160_1_42 = _q__idx_fsm___pip_5160_1_42;
_d__full_fsm___pip_5160_1_42 = _q__full_fsm___pip_5160_1_42;
_t__stall_fsm___pip_5160_1_42 = 0;
_t__1stdisable_fsm___pip_5160_1_42 = 0;
_d__idx_fsm___pip_5160_1_43 = _q__idx_fsm___pip_5160_1_43;
_d__full_fsm___pip_5160_1_43 = _q__full_fsm___pip_5160_1_43;
_t__stall_fsm___pip_5160_1_43 = 0;
_t__1stdisable_fsm___pip_5160_1_43 = 0;
_d__idx_fsm___pip_5160_1_44 = _q__idx_fsm___pip_5160_1_44;
_d__full_fsm___pip_5160_1_44 = _q__full_fsm___pip_5160_1_44;
_t__stall_fsm___pip_5160_1_44 = 0;
_t__1stdisable_fsm___pip_5160_1_44 = 0;
_d__idx_fsm___pip_5160_1_45 = _q__idx_fsm___pip_5160_1_45;
_d__full_fsm___pip_5160_1_45 = _q__full_fsm___pip_5160_1_45;
_t__stall_fsm___pip_5160_1_45 = 0;
_t__1stdisable_fsm___pip_5160_1_45 = 0;
_d__idx_fsm___pip_5160_1_46 = _q__idx_fsm___pip_5160_1_46;
_d__full_fsm___pip_5160_1_46 = _q__full_fsm___pip_5160_1_46;
_t__stall_fsm___pip_5160_1_46 = 0;
_t__1stdisable_fsm___pip_5160_1_46 = 0;
_d__idx_fsm___pip_5160_1_47 = _q__idx_fsm___pip_5160_1_47;
_d__full_fsm___pip_5160_1_47 = _q__full_fsm___pip_5160_1_47;
_t__stall_fsm___pip_5160_1_47 = 0;
_t__1stdisable_fsm___pip_5160_1_47 = 0;
_d__idx_fsm___pip_5160_1_48 = _q__idx_fsm___pip_5160_1_48;
_d__full_fsm___pip_5160_1_48 = _q__full_fsm___pip_5160_1_48;
_t__stall_fsm___pip_5160_1_48 = 0;
_t__1stdisable_fsm___pip_5160_1_48 = 0;
_d__idx_fsm___pip_5160_1_49 = _q__idx_fsm___pip_5160_1_49;
_d__full_fsm___pip_5160_1_49 = _q__full_fsm___pip_5160_1_49;
_t__stall_fsm___pip_5160_1_49 = 0;
_t__1stdisable_fsm___pip_5160_1_49 = 0;
_d__idx_fsm___pip_5160_1_50 = _q__idx_fsm___pip_5160_1_50;
_d__full_fsm___pip_5160_1_50 = _q__full_fsm___pip_5160_1_50;
_t__stall_fsm___pip_5160_1_50 = 0;
_t__1stdisable_fsm___pip_5160_1_50 = 0;
_d__idx_fsm___pip_5160_1_51 = _q__idx_fsm___pip_5160_1_51;
_d__full_fsm___pip_5160_1_51 = _q__full_fsm___pip_5160_1_51;
_t__stall_fsm___pip_5160_1_51 = 0;
_t__1stdisable_fsm___pip_5160_1_51 = 0;
_d__idx_fsm___pip_5160_1_52 = _q__idx_fsm___pip_5160_1_52;
_d__full_fsm___pip_5160_1_52 = _q__full_fsm___pip_5160_1_52;
_t__stall_fsm___pip_5160_1_52 = 0;
_t__1stdisable_fsm___pip_5160_1_52 = 0;
_d__idx_fsm___pip_5160_1_53 = _q__idx_fsm___pip_5160_1_53;
_d__full_fsm___pip_5160_1_53 = _q__full_fsm___pip_5160_1_53;
_t__stall_fsm___pip_5160_1_53 = 0;
_t__1stdisable_fsm___pip_5160_1_53 = 0;
_d__idx_fsm___pip_5160_1_54 = _q__idx_fsm___pip_5160_1_54;
_d__full_fsm___pip_5160_1_54 = _q__full_fsm___pip_5160_1_54;
_t__stall_fsm___pip_5160_1_54 = 0;
_t__1stdisable_fsm___pip_5160_1_54 = 0;
_d__idx_fsm___pip_5160_1_55 = _q__idx_fsm___pip_5160_1_55;
_d__full_fsm___pip_5160_1_55 = _q__full_fsm___pip_5160_1_55;
_t__stall_fsm___pip_5160_1_55 = 0;
_t__1stdisable_fsm___pip_5160_1_55 = 0;
_d__idx_fsm___pip_5160_1_56 = _q__idx_fsm___pip_5160_1_56;
_d__full_fsm___pip_5160_1_56 = _q__full_fsm___pip_5160_1_56;
_t__stall_fsm___pip_5160_1_56 = 0;
_t__1stdisable_fsm___pip_5160_1_56 = 0;
_d__idx_fsm___pip_5160_1_57 = _q__idx_fsm___pip_5160_1_57;
_d__full_fsm___pip_5160_1_57 = _q__full_fsm___pip_5160_1_57;
_t__stall_fsm___pip_5160_1_57 = 0;
_t__1stdisable_fsm___pip_5160_1_57 = 0;
_d__idx_fsm___pip_5160_1_58 = _q__idx_fsm___pip_5160_1_58;
_d__full_fsm___pip_5160_1_58 = _q__full_fsm___pip_5160_1_58;
_t__stall_fsm___pip_5160_1_58 = 0;
_t__1stdisable_fsm___pip_5160_1_58 = 0;
_d__idx_fsm___pip_5160_1_59 = _q__idx_fsm___pip_5160_1_59;
_d__full_fsm___pip_5160_1_59 = _q__full_fsm___pip_5160_1_59;
_t__stall_fsm___pip_5160_1_59 = 0;
_t__1stdisable_fsm___pip_5160_1_59 = 0;
_d__idx_fsm___pip_5160_1_60 = _q__idx_fsm___pip_5160_1_60;
_d__full_fsm___pip_5160_1_60 = _q__full_fsm___pip_5160_1_60;
_t__stall_fsm___pip_5160_1_60 = 0;
_t__1stdisable_fsm___pip_5160_1_60 = 0;
_d__idx_fsm___pip_5160_1_61 = _q__idx_fsm___pip_5160_1_61;
_d__full_fsm___pip_5160_1_61 = _q__full_fsm___pip_5160_1_61;
_t__stall_fsm___pip_5160_1_61 = 0;
_t__1stdisable_fsm___pip_5160_1_61 = 0;
_d__idx_fsm___pip_5160_1_62 = _q__idx_fsm___pip_5160_1_62;
_d__full_fsm___pip_5160_1_62 = _q__full_fsm___pip_5160_1_62;
_t__stall_fsm___pip_5160_1_62 = 0;
_t__1stdisable_fsm___pip_5160_1_62 = 0;
_d__idx_fsm___pip_5160_1_63 = _q__idx_fsm___pip_5160_1_63;
_d__full_fsm___pip_5160_1_63 = _q__full_fsm___pip_5160_1_63;
_t__stall_fsm___pip_5160_1_63 = 0;
_t__1stdisable_fsm___pip_5160_1_63 = 0;
_d__idx_fsm___pip_5160_1_64 = _q__idx_fsm___pip_5160_1_64;
_d__full_fsm___pip_5160_1_64 = _q__full_fsm___pip_5160_1_64;
_t__stall_fsm___pip_5160_1_64 = 0;
_t__1stdisable_fsm___pip_5160_1_64 = 0;
_d__idx_fsm___pip_5160_1_65 = _q__idx_fsm___pip_5160_1_65;
_d__full_fsm___pip_5160_1_65 = _q__full_fsm___pip_5160_1_65;
_t__stall_fsm___pip_5160_1_65 = 0;
_t__1stdisable_fsm___pip_5160_1_65 = 0;
_d__idx_fsm___pip_5160_1_66 = _q__idx_fsm___pip_5160_1_66;
_d__full_fsm___pip_5160_1_66 = _q__full_fsm___pip_5160_1_66;
_t__stall_fsm___pip_5160_1_66 = 0;
_t__1stdisable_fsm___pip_5160_1_66 = 0;
_d__idx_fsm___pip_5160_1_67 = _q__idx_fsm___pip_5160_1_67;
_d__full_fsm___pip_5160_1_67 = _q__full_fsm___pip_5160_1_67;
_t__stall_fsm___pip_5160_1_67 = 0;
_t__1stdisable_fsm___pip_5160_1_67 = 0;
_d__idx_fsm___pip_5160_1_68 = _q__idx_fsm___pip_5160_1_68;
_d__full_fsm___pip_5160_1_68 = _q__full_fsm___pip_5160_1_68;
_t__stall_fsm___pip_5160_1_68 = 0;
_t__1stdisable_fsm___pip_5160_1_68 = 0;
_d__idx_fsm___pip_5160_1_69 = _q__idx_fsm___pip_5160_1_69;
_d__full_fsm___pip_5160_1_69 = _q__full_fsm___pip_5160_1_69;
_t__stall_fsm___pip_5160_1_69 = 0;
_t__1stdisable_fsm___pip_5160_1_69 = 0;
_d__idx_fsm___pip_5160_1_70 = _q__idx_fsm___pip_5160_1_70;
_d__full_fsm___pip_5160_1_70 = _q__full_fsm___pip_5160_1_70;
_t__stall_fsm___pip_5160_1_70 = 0;
_t__1stdisable_fsm___pip_5160_1_70 = 0;
_d__idx_fsm___pip_5160_1_71 = _q__idx_fsm___pip_5160_1_71;
_d__full_fsm___pip_5160_1_71 = _q__full_fsm___pip_5160_1_71;
_t__stall_fsm___pip_5160_1_71 = 0;
_t__1stdisable_fsm___pip_5160_1_71 = 0;
_d__idx_fsm___pip_5160_1_72 = _q__idx_fsm___pip_5160_1_72;
_d__full_fsm___pip_5160_1_72 = _q__full_fsm___pip_5160_1_72;
_t__stall_fsm___pip_5160_1_72 = 0;
_t__1stdisable_fsm___pip_5160_1_72 = 0;
_d__idx_fsm___pip_5160_1_73 = _q__idx_fsm___pip_5160_1_73;
_d__full_fsm___pip_5160_1_73 = _q__full_fsm___pip_5160_1_73;
_t__stall_fsm___pip_5160_1_73 = 0;
_t__1stdisable_fsm___pip_5160_1_73 = 0;
_d__idx_fsm___pip_5160_1_74 = _q__idx_fsm___pip_5160_1_74;
_d__full_fsm___pip_5160_1_74 = _q__full_fsm___pip_5160_1_74;
_t__stall_fsm___pip_5160_1_74 = 0;
_t__1stdisable_fsm___pip_5160_1_74 = 0;
_d__idx_fsm___pip_5160_1_75 = _q__idx_fsm___pip_5160_1_75;
_d__full_fsm___pip_5160_1_75 = _q__full_fsm___pip_5160_1_75;
_t__stall_fsm___pip_5160_1_75 = 0;
_t__1stdisable_fsm___pip_5160_1_75 = 0;
_d__idx_fsm___pip_5160_1_76 = _q__idx_fsm___pip_5160_1_76;
_d__full_fsm___pip_5160_1_76 = _q__full_fsm___pip_5160_1_76;
_t__stall_fsm___pip_5160_1_76 = 0;
_t__1stdisable_fsm___pip_5160_1_76 = 0;
_d__idx_fsm___pip_5160_1_77 = _q__idx_fsm___pip_5160_1_77;
_d__full_fsm___pip_5160_1_77 = _q__full_fsm___pip_5160_1_77;
_t__stall_fsm___pip_5160_1_77 = 0;
_t__1stdisable_fsm___pip_5160_1_77 = 0;
_d__idx_fsm___pip_5160_1_78 = _q__idx_fsm___pip_5160_1_78;
_d__full_fsm___pip_5160_1_78 = _q__full_fsm___pip_5160_1_78;
_t__stall_fsm___pip_5160_1_78 = 0;
_t__1stdisable_fsm___pip_5160_1_78 = 0;
_d__idx_fsm___pip_5160_1_79 = _q__idx_fsm___pip_5160_1_79;
_d__full_fsm___pip_5160_1_79 = _q__full_fsm___pip_5160_1_79;
_t__stall_fsm___pip_5160_1_79 = 0;
_t__1stdisable_fsm___pip_5160_1_79 = 0;
_d__idx_fsm___pip_5160_1_80 = _q__idx_fsm___pip_5160_1_80;
_d__full_fsm___pip_5160_1_80 = _q__full_fsm___pip_5160_1_80;
_t__stall_fsm___pip_5160_1_80 = 0;
_t__1stdisable_fsm___pip_5160_1_80 = 0;
_d__idx_fsm___pip_5160_1_81 = _q__idx_fsm___pip_5160_1_81;
_d__full_fsm___pip_5160_1_81 = _q__full_fsm___pip_5160_1_81;
_t__stall_fsm___pip_5160_1_81 = 0;
_t__1stdisable_fsm___pip_5160_1_81 = 0;
_d__idx_fsm___pip_5160_1_82 = _q__idx_fsm___pip_5160_1_82;
_d__full_fsm___pip_5160_1_82 = _q__full_fsm___pip_5160_1_82;
_t__stall_fsm___pip_5160_1_82 = 0;
_t__1stdisable_fsm___pip_5160_1_82 = 0;
_d__idx_fsm___pip_5160_1_83 = _q__idx_fsm___pip_5160_1_83;
_d__full_fsm___pip_5160_1_83 = _q__full_fsm___pip_5160_1_83;
_t__stall_fsm___pip_5160_1_83 = 0;
_t__1stdisable_fsm___pip_5160_1_83 = 0;
_d__idx_fsm___pip_5160_1_84 = _q__idx_fsm___pip_5160_1_84;
_d__full_fsm___pip_5160_1_84 = _q__full_fsm___pip_5160_1_84;
_t__stall_fsm___pip_5160_1_84 = 0;
_t__1stdisable_fsm___pip_5160_1_84 = 0;
_d__idx_fsm___pip_5160_1_85 = _q__idx_fsm___pip_5160_1_85;
_d__full_fsm___pip_5160_1_85 = _q__full_fsm___pip_5160_1_85;
_t__stall_fsm___pip_5160_1_85 = 0;
_t__1stdisable_fsm___pip_5160_1_85 = 0;
_d__idx_fsm___pip_5160_1_86 = _q__idx_fsm___pip_5160_1_86;
_d__full_fsm___pip_5160_1_86 = _q__full_fsm___pip_5160_1_86;
_t__stall_fsm___pip_5160_1_86 = 0;
_t__1stdisable_fsm___pip_5160_1_86 = 0;
_d__idx_fsm___pip_5160_1_87 = _q__idx_fsm___pip_5160_1_87;
_d__full_fsm___pip_5160_1_87 = _q__full_fsm___pip_5160_1_87;
_t__stall_fsm___pip_5160_1_87 = 0;
_t__1stdisable_fsm___pip_5160_1_87 = 0;
_d__idx_fsm___pip_5160_1_88 = _q__idx_fsm___pip_5160_1_88;
_d__full_fsm___pip_5160_1_88 = _q__full_fsm___pip_5160_1_88;
_t__stall_fsm___pip_5160_1_88 = 0;
_t__1stdisable_fsm___pip_5160_1_88 = 0;
_d__idx_fsm___pip_5160_1_89 = _q__idx_fsm___pip_5160_1_89;
_d__full_fsm___pip_5160_1_89 = _q__full_fsm___pip_5160_1_89;
_t__stall_fsm___pip_5160_1_89 = 0;
_t__1stdisable_fsm___pip_5160_1_89 = 0;
_d__idx_fsm___pip_5160_1_90 = _q__idx_fsm___pip_5160_1_90;
_d__full_fsm___pip_5160_1_90 = _q__full_fsm___pip_5160_1_90;
_t__stall_fsm___pip_5160_1_90 = 0;
_t__1stdisable_fsm___pip_5160_1_90 = 0;
_d__idx_fsm___pip_5160_1_91 = _q__idx_fsm___pip_5160_1_91;
_d__full_fsm___pip_5160_1_91 = _q__full_fsm___pip_5160_1_91;
_t__stall_fsm___pip_5160_1_91 = 0;
_t__1stdisable_fsm___pip_5160_1_91 = 0;
_d__idx_fsm___pip_5160_1_92 = _q__idx_fsm___pip_5160_1_92;
_d__full_fsm___pip_5160_1_92 = _q__full_fsm___pip_5160_1_92;
_t__stall_fsm___pip_5160_1_92 = 0;
_t__1stdisable_fsm___pip_5160_1_92 = 0;
_d__idx_fsm___pip_5160_1_93 = _q__idx_fsm___pip_5160_1_93;
_d__full_fsm___pip_5160_1_93 = _q__full_fsm___pip_5160_1_93;
_t__stall_fsm___pip_5160_1_93 = 0;
_t__1stdisable_fsm___pip_5160_1_93 = 0;
_d__idx_fsm___pip_5160_1_94 = _q__idx_fsm___pip_5160_1_94;
_d__full_fsm___pip_5160_1_94 = _q__full_fsm___pip_5160_1_94;
_t__stall_fsm___pip_5160_1_94 = 0;
_t__1stdisable_fsm___pip_5160_1_94 = 0;
_d__idx_fsm___pip_5160_1_95 = _q__idx_fsm___pip_5160_1_95;
_d__full_fsm___pip_5160_1_95 = _q__full_fsm___pip_5160_1_95;
_t__stall_fsm___pip_5160_1_95 = 0;
_t__1stdisable_fsm___pip_5160_1_95 = 0;
_d__idx_fsm___pip_5160_1_96 = _q__idx_fsm___pip_5160_1_96;
_d__full_fsm___pip_5160_1_96 = _q__full_fsm___pip_5160_1_96;
_t__stall_fsm___pip_5160_1_96 = 0;
_t__1stdisable_fsm___pip_5160_1_96 = 0;
_d__idx_fsm___pip_5160_1_97 = _q__idx_fsm___pip_5160_1_97;
_d__full_fsm___pip_5160_1_97 = _q__full_fsm___pip_5160_1_97;
_t__stall_fsm___pip_5160_1_97 = 0;
_t__1stdisable_fsm___pip_5160_1_97 = 0;
_d__idx_fsm___pip_5160_1_98 = _q__idx_fsm___pip_5160_1_98;
_d__full_fsm___pip_5160_1_98 = _q__full_fsm___pip_5160_1_98;
_t__stall_fsm___pip_5160_1_98 = 0;
_t__1stdisable_fsm___pip_5160_1_98 = 0;
_d__idx_fsm___pip_5160_1_99 = _q__idx_fsm___pip_5160_1_99;
_d__full_fsm___pip_5160_1_99 = _q__full_fsm___pip_5160_1_99;
_t__stall_fsm___pip_5160_1_99 = 0;
_t__1stdisable_fsm___pip_5160_1_99 = 0;
_d__idx_fsm___pip_5160_1_100 = _q__idx_fsm___pip_5160_1_100;
_d__full_fsm___pip_5160_1_100 = _q__full_fsm___pip_5160_1_100;
_t__stall_fsm___pip_5160_1_100 = 0;
_t__1stdisable_fsm___pip_5160_1_100 = 0;
_d__idx_fsm___pip_5160_1_101 = _q__idx_fsm___pip_5160_1_101;
_d__full_fsm___pip_5160_1_101 = _q__full_fsm___pip_5160_1_101;
_t__stall_fsm___pip_5160_1_101 = 0;
_t__1stdisable_fsm___pip_5160_1_101 = 0;
_d__idx_fsm___pip_5160_1_102 = _q__idx_fsm___pip_5160_1_102;
_d__full_fsm___pip_5160_1_102 = _q__full_fsm___pip_5160_1_102;
_t__stall_fsm___pip_5160_1_102 = 0;
_t__1stdisable_fsm___pip_5160_1_102 = 0;
_d__idx_fsm___pip_5160_1_103 = _q__idx_fsm___pip_5160_1_103;
_d__full_fsm___pip_5160_1_103 = _q__full_fsm___pip_5160_1_103;
_t__stall_fsm___pip_5160_1_103 = 0;
_t__1stdisable_fsm___pip_5160_1_103 = 0;
_d__idx_fsm___pip_5160_1_104 = _q__idx_fsm___pip_5160_1_104;
_d__full_fsm___pip_5160_1_104 = _q__full_fsm___pip_5160_1_104;
_t__stall_fsm___pip_5160_1_104 = 0;
_t__1stdisable_fsm___pip_5160_1_104 = 0;
_d__idx_fsm___pip_5160_1_105 = _q__idx_fsm___pip_5160_1_105;
_d__full_fsm___pip_5160_1_105 = _q__full_fsm___pip_5160_1_105;
_t__stall_fsm___pip_5160_1_105 = 0;
_t__1stdisable_fsm___pip_5160_1_105 = 0;
_d__idx_fsm___pip_5160_1_106 = _q__idx_fsm___pip_5160_1_106;
_d__full_fsm___pip_5160_1_106 = _q__full_fsm___pip_5160_1_106;
_t__stall_fsm___pip_5160_1_106 = 0;
_t__1stdisable_fsm___pip_5160_1_106 = 0;
_d__idx_fsm___pip_5160_1_107 = _q__idx_fsm___pip_5160_1_107;
_d__full_fsm___pip_5160_1_107 = _q__full_fsm___pip_5160_1_107;
_t__stall_fsm___pip_5160_1_107 = 0;
_t__1stdisable_fsm___pip_5160_1_107 = 0;
_d__idx_fsm___pip_5160_1_108 = _q__idx_fsm___pip_5160_1_108;
_d__full_fsm___pip_5160_1_108 = _q__full_fsm___pip_5160_1_108;
_t__stall_fsm___pip_5160_1_108 = 0;
_t__1stdisable_fsm___pip_5160_1_108 = 0;
_d__idx_fsm___pip_5160_1_109 = _q__idx_fsm___pip_5160_1_109;
_d__full_fsm___pip_5160_1_109 = _q__full_fsm___pip_5160_1_109;
_t__stall_fsm___pip_5160_1_109 = 0;
_t__1stdisable_fsm___pip_5160_1_109 = 0;
_d__idx_fsm___pip_5160_1_110 = _q__idx_fsm___pip_5160_1_110;
_d__full_fsm___pip_5160_1_110 = _q__full_fsm___pip_5160_1_110;
_t__stall_fsm___pip_5160_1_110 = 0;
_t__1stdisable_fsm___pip_5160_1_110 = 0;
_d__idx_fsm___pip_5160_1_111 = _q__idx_fsm___pip_5160_1_111;
_d__full_fsm___pip_5160_1_111 = _q__full_fsm___pip_5160_1_111;
_t__stall_fsm___pip_5160_1_111 = 0;
_t__1stdisable_fsm___pip_5160_1_111 = 0;
_d__idx_fsm___pip_5160_1_112 = _q__idx_fsm___pip_5160_1_112;
_d__full_fsm___pip_5160_1_112 = _q__full_fsm___pip_5160_1_112;
_t__stall_fsm___pip_5160_1_112 = 0;
_t__1stdisable_fsm___pip_5160_1_112 = 0;
_d__idx_fsm___pip_5160_1_113 = _q__idx_fsm___pip_5160_1_113;
_d__full_fsm___pip_5160_1_113 = _q__full_fsm___pip_5160_1_113;
_t__stall_fsm___pip_5160_1_113 = 0;
_t__1stdisable_fsm___pip_5160_1_113 = 0;
_d__idx_fsm___pip_5160_1_114 = _q__idx_fsm___pip_5160_1_114;
_d__full_fsm___pip_5160_1_114 = _q__full_fsm___pip_5160_1_114;
_t__stall_fsm___pip_5160_1_114 = 0;
_t__1stdisable_fsm___pip_5160_1_114 = 0;
_d__idx_fsm___pip_5160_1_115 = _q__idx_fsm___pip_5160_1_115;
_d__full_fsm___pip_5160_1_115 = _q__full_fsm___pip_5160_1_115;
_t__stall_fsm___pip_5160_1_115 = 0;
_t__1stdisable_fsm___pip_5160_1_115 = 0;
_d__idx_fsm___pip_5160_1_116 = _q__idx_fsm___pip_5160_1_116;
_d__full_fsm___pip_5160_1_116 = _q__full_fsm___pip_5160_1_116;
_t__stall_fsm___pip_5160_1_116 = 0;
_t__1stdisable_fsm___pip_5160_1_116 = 0;
_d__idx_fsm___pip_5160_1_117 = _q__idx_fsm___pip_5160_1_117;
_d__full_fsm___pip_5160_1_117 = _q__full_fsm___pip_5160_1_117;
_t__stall_fsm___pip_5160_1_117 = 0;
_t__1stdisable_fsm___pip_5160_1_117 = 0;
_d__idx_fsm___pip_5160_1_118 = _q__idx_fsm___pip_5160_1_118;
_d__full_fsm___pip_5160_1_118 = _q__full_fsm___pip_5160_1_118;
_t__stall_fsm___pip_5160_1_118 = 0;
_t__1stdisable_fsm___pip_5160_1_118 = 0;
_d__idx_fsm___pip_5160_1_119 = _q__idx_fsm___pip_5160_1_119;
_d__full_fsm___pip_5160_1_119 = _q__full_fsm___pip_5160_1_119;
_t__stall_fsm___pip_5160_1_119 = 0;
_t__1stdisable_fsm___pip_5160_1_119 = 0;
_d__idx_fsm___pip_5160_1_120 = _q__idx_fsm___pip_5160_1_120;
_d__full_fsm___pip_5160_1_120 = _q__full_fsm___pip_5160_1_120;
_t__stall_fsm___pip_5160_1_120 = 0;
_t__1stdisable_fsm___pip_5160_1_120 = 0;
_d__idx_fsm___pip_5160_1_121 = _q__idx_fsm___pip_5160_1_121;
_d__full_fsm___pip_5160_1_121 = _q__full_fsm___pip_5160_1_121;
_t__stall_fsm___pip_5160_1_121 = 0;
_t__1stdisable_fsm___pip_5160_1_121 = 0;
_d__idx_fsm___pip_5160_1_122 = _q__idx_fsm___pip_5160_1_122;
_d__full_fsm___pip_5160_1_122 = _q__full_fsm___pip_5160_1_122;
_t__stall_fsm___pip_5160_1_122 = 0;
_t__1stdisable_fsm___pip_5160_1_122 = 0;
_d__idx_fsm___pip_5160_1_123 = _q__idx_fsm___pip_5160_1_123;
_d__full_fsm___pip_5160_1_123 = _q__full_fsm___pip_5160_1_123;
_t__stall_fsm___pip_5160_1_123 = 0;
_t__1stdisable_fsm___pip_5160_1_123 = 0;
_d__idx_fsm___pip_5160_1_124 = _q__idx_fsm___pip_5160_1_124;
_d__full_fsm___pip_5160_1_124 = _q__full_fsm___pip_5160_1_124;
_t__stall_fsm___pip_5160_1_124 = 0;
_t__1stdisable_fsm___pip_5160_1_124 = 0;
_d__idx_fsm___pip_5160_1_125 = _q__idx_fsm___pip_5160_1_125;
_d__full_fsm___pip_5160_1_125 = _q__full_fsm___pip_5160_1_125;
_t__stall_fsm___pip_5160_1_125 = 0;
_t__1stdisable_fsm___pip_5160_1_125 = 0;
_d__idx_fsm___pip_5160_1_126 = _q__idx_fsm___pip_5160_1_126;
_d__full_fsm___pip_5160_1_126 = _q__full_fsm___pip_5160_1_126;
_t__stall_fsm___pip_5160_1_126 = 0;
_t__1stdisable_fsm___pip_5160_1_126 = 0;
_d__idx_fsm___pip_5160_1_127 = _q__idx_fsm___pip_5160_1_127;
_d__full_fsm___pip_5160_1_127 = _q__full_fsm___pip_5160_1_127;
_t__stall_fsm___pip_5160_1_127 = 0;
_t__1stdisable_fsm___pip_5160_1_127 = 0;
_d__idx_fsm___pip_5160_1_128 = _q__idx_fsm___pip_5160_1_128;
_d__full_fsm___pip_5160_1_128 = _q__full_fsm___pip_5160_1_128;
_t__stall_fsm___pip_5160_1_128 = 0;
_t__1stdisable_fsm___pip_5160_1_128 = 0;
_d__idx_fsm___pip_5160_1_129 = _q__idx_fsm___pip_5160_1_129;
_d__full_fsm___pip_5160_1_129 = _q__full_fsm___pip_5160_1_129;
_t__stall_fsm___pip_5160_1_129 = 0;
_t__1stdisable_fsm___pip_5160_1_129 = 0;
_d__idx_fsm___pip_5160_1_130 = _q__idx_fsm___pip_5160_1_130;
_d__full_fsm___pip_5160_1_130 = _q__full_fsm___pip_5160_1_130;
_t__stall_fsm___pip_5160_1_130 = 0;
_t__1stdisable_fsm___pip_5160_1_130 = 0;
_d__idx_fsm___pip_5160_1_131 = _q__idx_fsm___pip_5160_1_131;
_d__full_fsm___pip_5160_1_131 = _q__full_fsm___pip_5160_1_131;
_t__stall_fsm___pip_5160_1_131 = 0;
_t__1stdisable_fsm___pip_5160_1_131 = 0;
_d__idx_fsm___pip_5160_1_132 = _q__idx_fsm___pip_5160_1_132;
_d__full_fsm___pip_5160_1_132 = _q__full_fsm___pip_5160_1_132;
_t__stall_fsm___pip_5160_1_132 = 0;
_t__1stdisable_fsm___pip_5160_1_132 = 0;
_d__idx_fsm___pip_5160_1_133 = _q__idx_fsm___pip_5160_1_133;
_d__full_fsm___pip_5160_1_133 = _q__full_fsm___pip_5160_1_133;
_t__stall_fsm___pip_5160_1_133 = 0;
_t__1stdisable_fsm___pip_5160_1_133 = 0;
_d__idx_fsm___pip_5160_1_134 = _q__idx_fsm___pip_5160_1_134;
_d__full_fsm___pip_5160_1_134 = _q__full_fsm___pip_5160_1_134;
_t__stall_fsm___pip_5160_1_134 = 0;
_t__1stdisable_fsm___pip_5160_1_134 = 0;
_d__idx_fsm___pip_5160_1_135 = _q__idx_fsm___pip_5160_1_135;
_d__full_fsm___pip_5160_1_135 = _q__full_fsm___pip_5160_1_135;
_t__stall_fsm___pip_5160_1_135 = 0;
_t__1stdisable_fsm___pip_5160_1_135 = 0;
_d__idx_fsm___pip_5160_1_136 = _q__idx_fsm___pip_5160_1_136;
_d__full_fsm___pip_5160_1_136 = _q__full_fsm___pip_5160_1_136;
_t__stall_fsm___pip_5160_1_136 = 0;
_t__1stdisable_fsm___pip_5160_1_136 = 0;
_t_cos_wenable0 = 0;
_t_cos_wdata0 = 0;
_t_cos_wenable1 = 0;
_t_cos_wdata1 = 0;
_t_sin_wenable0 = 0;
_t_sin_wdata0 = 0;
_t_sin_wenable1 = 0;
_t_sin_wdata1 = 0;
_t_invA_wenable0 = 0;
_t_invA_wdata0 = 0;
_t_invA_wenable1 = 0;
_t_invA_wdata1 = 0;
_t_invB_wenable = 0;
_t_invB_wdata = 0;
_t___stage___block_6_vxsz = 0;
_t___stage___block_6_view_x = 0;
_t___stage___block_6_view_y = 0;
_t___stage___block_7_cs0 = 0;
_t___stage___block_7_ss0 = 0;
_t___stage___block_7_cs1 = 0;
_t___stage___block_7_ss1 = 0;
_t___stage___block_7_rot_x = 0;
_t___stage___block_7_rot_y = 0;
_t___block_11_ycs = 0;
_t___block_11_yss = 0;
_t___stage___block_17_xcs = 0;
_t___block_19_xss = 0;
_t___block_21_zcs = 0;
_t___block_23_zss = 0;
_t___block_25_r_x_delta = 0;
_t___block_25_r_z_delta = 0;
_t___stage___block_26_rd_x = 0;
_t___stage___block_26_rd_y = 0;
_t___stage___block_26_rd_z = 0;
_t___stage___block_26_s_x = 0;
_t___stage___block_26_s_y = 0;
_t___stage___block_26_s_z = 0;
_t___stage___block_26_p_x = 0;
_t___stage___block_26_p_y = 0;
_t___stage___block_26_p_z = 0;
_t___stage___block_26_v_x = 0;
_t___stage___block_26_v_y = 0;
_t___stage___block_26_v_z = 0;
_t___stage___block_26_brd_x = 0;
_t___stage___block_26_brd_y = 0;
_t___stage___block_26_brd_z = 0;
_t___stage___block_28_inv_x = 0;
_t___stage___block_28_inv_y = 0;
_t___stage___block_28_inv_z = 0;
_t___stage___block_28_tm_x_ = 0;
_t___stage___block_28_tm_y_ = 0;
_t___stage___block_28_tm_z_ = 0;
_t___block_34_tm_x = 0;
_t___block_34_tm_y = 0;
_t___block_34_tm_z = 0;
_t___block_34_dt_x_ = 0;
_t___block_34_dt_y_ = 0;
_t___block_34_dt_z_ = 0;
_t___block_40_dt_x = 0;
_t___block_40_dt_y = 0;
_t___block_40_dt_z = 0;
_t___stage___block_41_tex = 0;
_t___stage___block_41_vnum0 = 0;
_t___stage___block_41_vnum1 = 0;
_t___stage___block_41_vnum2 = 0;
_t___block_46_cmp_yx = 0;
_t___block_46_cmp_zx = 0;
_t___block_46_cmp_zy = 0;
_t___block_46_x_sel = 0;
_t___block_46_y_sel = 0;
_t___block_46_z_sel = 0;
_t___stage___block_62_tex = 0;
_t___stage___block_62_vnum0 = 0;
_t___stage___block_62_vnum1 = 0;
_t___stage___block_62_vnum2 = 0;
_t___block_67_cmp_yx = 0;
_t___block_67_cmp_zx = 0;
_t___block_67_cmp_zy = 0;
_t___block_67_x_sel = 0;
_t___block_67_y_sel = 0;
_t___block_67_z_sel = 0;
_t___stage___block_83_tex = 0;
_t___stage___block_83_vnum0 = 0;
_t___stage___block_83_vnum1 = 0;
_t___stage___block_83_vnum2 = 0;
_t___block_88_cmp_yx = 0;
_t___block_88_cmp_zx = 0;
_t___block_88_cmp_zy = 0;
_t___block_88_x_sel = 0;
_t___block_88_y_sel = 0;
_t___block_88_z_sel = 0;
_t___stage___block_104_tex = 0;
_t___stage___block_104_vnum0 = 0;
_t___stage___block_104_vnum1 = 0;
_t___stage___block_104_vnum2 = 0;
_t___block_109_cmp_yx = 0;
_t___block_109_cmp_zx = 0;
_t___block_109_cmp_zy = 0;
_t___block_109_x_sel = 0;
_t___block_109_y_sel = 0;
_t___block_109_z_sel = 0;
_t___stage___block_125_tex = 0;
_t___stage___block_125_vnum0 = 0;
_t___stage___block_125_vnum1 = 0;
_t___stage___block_125_vnum2 = 0;
_t___block_130_cmp_yx = 0;
_t___block_130_cmp_zx = 0;
_t___block_130_cmp_zy = 0;
_t___block_130_x_sel = 0;
_t___block_130_y_sel = 0;
_t___block_130_z_sel = 0;
_t___stage___block_146_tex = 0;
_t___stage___block_146_vnum0 = 0;
_t___stage___block_146_vnum1 = 0;
_t___stage___block_146_vnum2 = 0;
_t___block_151_cmp_yx = 0;
_t___block_151_cmp_zx = 0;
_t___block_151_cmp_zy = 0;
_t___block_151_x_sel = 0;
_t___block_151_y_sel = 0;
_t___block_151_z_sel = 0;
_t___stage___block_167_tex = 0;
_t___stage___block_167_vnum0 = 0;
_t___stage___block_167_vnum1 = 0;
_t___stage___block_167_vnum2 = 0;
_t___block_172_cmp_yx = 0;
_t___block_172_cmp_zx = 0;
_t___block_172_cmp_zy = 0;
_t___block_172_x_sel = 0;
_t___block_172_y_sel = 0;
_t___block_172_z_sel = 0;
_t___stage___block_188_tex = 0;
_t___stage___block_188_vnum0 = 0;
_t___stage___block_188_vnum1 = 0;
_t___stage___block_188_vnum2 = 0;
_t___block_193_cmp_yx = 0;
_t___block_193_cmp_zx = 0;
_t___block_193_cmp_zy = 0;
_t___block_193_x_sel = 0;
_t___block_193_y_sel = 0;
_t___block_193_z_sel = 0;
_t___stage___block_209_tex = 0;
_t___stage___block_209_vnum0 = 0;
_t___stage___block_209_vnum1 = 0;
_t___stage___block_209_vnum2 = 0;
_t___block_214_cmp_yx = 0;
_t___block_214_cmp_zx = 0;
_t___block_214_cmp_zy = 0;
_t___block_214_x_sel = 0;
_t___block_214_y_sel = 0;
_t___block_214_z_sel = 0;
_t___stage___block_230_tex = 0;
_t___stage___block_230_vnum0 = 0;
_t___stage___block_230_vnum1 = 0;
_t___stage___block_230_vnum2 = 0;
_t___block_235_cmp_yx = 0;
_t___block_235_cmp_zx = 0;
_t___block_235_cmp_zy = 0;
_t___block_235_x_sel = 0;
_t___block_235_y_sel = 0;
_t___block_235_z_sel = 0;
_t___stage___block_251_tex = 0;
_t___stage___block_251_vnum0 = 0;
_t___stage___block_251_vnum1 = 0;
_t___stage___block_251_vnum2 = 0;
_t___block_256_cmp_yx = 0;
_t___block_256_cmp_zx = 0;
_t___block_256_cmp_zy = 0;
_t___block_256_x_sel = 0;
_t___block_256_y_sel = 0;
_t___block_256_z_sel = 0;
_t___stage___block_272_tex = 0;
_t___stage___block_272_vnum0 = 0;
_t___stage___block_272_vnum1 = 0;
_t___stage___block_272_vnum2 = 0;
_t___block_277_cmp_yx = 0;
_t___block_277_cmp_zx = 0;
_t___block_277_cmp_zy = 0;
_t___block_277_x_sel = 0;
_t___block_277_y_sel = 0;
_t___block_277_z_sel = 0;
_t___stage___block_293_tex = 0;
_t___stage___block_293_vnum0 = 0;
_t___stage___block_293_vnum1 = 0;
_t___stage___block_293_vnum2 = 0;
_t___block_298_cmp_yx = 0;
_t___block_298_cmp_zx = 0;
_t___block_298_cmp_zy = 0;
_t___block_298_x_sel = 0;
_t___block_298_y_sel = 0;
_t___block_298_z_sel = 0;
_t___stage___block_314_tex = 0;
_t___stage___block_314_vnum0 = 0;
_t___stage___block_314_vnum1 = 0;
_t___stage___block_314_vnum2 = 0;
_t___block_319_cmp_yx = 0;
_t___block_319_cmp_zx = 0;
_t___block_319_cmp_zy = 0;
_t___block_319_x_sel = 0;
_t___block_319_y_sel = 0;
_t___block_319_z_sel = 0;
_t___stage___block_335_tex = 0;
_t___stage___block_335_vnum0 = 0;
_t___stage___block_335_vnum1 = 0;
_t___stage___block_335_vnum2 = 0;
_t___block_340_cmp_yx = 0;
_t___block_340_cmp_zx = 0;
_t___block_340_cmp_zy = 0;
_t___block_340_x_sel = 0;
_t___block_340_y_sel = 0;
_t___block_340_z_sel = 0;
_t___stage___block_356_tex = 0;
_t___stage___block_356_vnum0 = 0;
_t___stage___block_356_vnum1 = 0;
_t___stage___block_356_vnum2 = 0;
_t___block_361_cmp_yx = 0;
_t___block_361_cmp_zx = 0;
_t___block_361_cmp_zy = 0;
_t___block_361_x_sel = 0;
_t___block_361_y_sel = 0;
_t___block_361_z_sel = 0;
_t___stage___block_377_tex = 0;
_t___stage___block_377_vnum0 = 0;
_t___stage___block_377_vnum1 = 0;
_t___stage___block_377_vnum2 = 0;
_t___block_382_cmp_yx = 0;
_t___block_382_cmp_zx = 0;
_t___block_382_cmp_zy = 0;
_t___block_382_x_sel = 0;
_t___block_382_y_sel = 0;
_t___block_382_z_sel = 0;
_t___stage___block_398_tex = 0;
_t___stage___block_398_vnum0 = 0;
_t___stage___block_398_vnum1 = 0;
_t___stage___block_398_vnum2 = 0;
_t___block_403_cmp_yx = 0;
_t___block_403_cmp_zx = 0;
_t___block_403_cmp_zy = 0;
_t___block_403_x_sel = 0;
_t___block_403_y_sel = 0;
_t___block_403_z_sel = 0;
_t___stage___block_419_tex = 0;
_t___stage___block_419_vnum0 = 0;
_t___stage___block_419_vnum1 = 0;
_t___stage___block_419_vnum2 = 0;
_t___block_424_cmp_yx = 0;
_t___block_424_cmp_zx = 0;
_t___block_424_cmp_zy = 0;
_t___block_424_x_sel = 0;
_t___block_424_y_sel = 0;
_t___block_424_z_sel = 0;
_t___stage___block_440_tex = 0;
_t___stage___block_440_vnum0 = 0;
_t___stage___block_440_vnum1 = 0;
_t___stage___block_440_vnum2 = 0;
_t___block_445_cmp_yx = 0;
_t___block_445_cmp_zx = 0;
_t___block_445_cmp_zy = 0;
_t___block_445_x_sel = 0;
_t___block_445_y_sel = 0;
_t___block_445_z_sel = 0;
_t___stage___block_461_tex = 0;
_t___stage___block_461_vnum0 = 0;
_t___stage___block_461_vnum1 = 0;
_t___stage___block_461_vnum2 = 0;
_t___block_466_cmp_yx = 0;
_t___block_466_cmp_zx = 0;
_t___block_466_cmp_zy = 0;
_t___block_466_x_sel = 0;
_t___block_466_y_sel = 0;
_t___block_466_z_sel = 0;
_t___stage___block_482_tex = 0;
_t___stage___block_482_vnum0 = 0;
_t___stage___block_482_vnum1 = 0;
_t___stage___block_482_vnum2 = 0;
_t___block_487_cmp_yx = 0;
_t___block_487_cmp_zx = 0;
_t___block_487_cmp_zy = 0;
_t___block_487_x_sel = 0;
_t___block_487_y_sel = 0;
_t___block_487_z_sel = 0;
_t___stage___block_503_tex = 0;
_t___stage___block_503_vnum0 = 0;
_t___stage___block_503_vnum1 = 0;
_t___stage___block_503_vnum2 = 0;
_t___block_508_cmp_yx = 0;
_t___block_508_cmp_zx = 0;
_t___block_508_cmp_zy = 0;
_t___block_508_x_sel = 0;
_t___block_508_y_sel = 0;
_t___block_508_z_sel = 0;
_t___stage___block_524_tex = 0;
_t___stage___block_524_vnum0 = 0;
_t___stage___block_524_vnum1 = 0;
_t___stage___block_524_vnum2 = 0;
_t___block_529_cmp_yx = 0;
_t___block_529_cmp_zx = 0;
_t___block_529_cmp_zy = 0;
_t___block_529_x_sel = 0;
_t___block_529_y_sel = 0;
_t___block_529_z_sel = 0;
_t___stage___block_545_tex = 0;
_t___stage___block_545_vnum0 = 0;
_t___stage___block_545_vnum1 = 0;
_t___stage___block_545_vnum2 = 0;
_t___block_550_cmp_yx = 0;
_t___block_550_cmp_zx = 0;
_t___block_550_cmp_zy = 0;
_t___block_550_x_sel = 0;
_t___block_550_y_sel = 0;
_t___block_550_z_sel = 0;
_t___stage___block_566_tex = 0;
_t___stage___block_566_vnum0 = 0;
_t___stage___block_566_vnum1 = 0;
_t___stage___block_566_vnum2 = 0;
_t___block_571_cmp_yx = 0;
_t___block_571_cmp_zx = 0;
_t___block_571_cmp_zy = 0;
_t___block_571_x_sel = 0;
_t___block_571_y_sel = 0;
_t___block_571_z_sel = 0;
_t___stage___block_587_tex = 0;
_t___stage___block_587_vnum0 = 0;
_t___stage___block_587_vnum1 = 0;
_t___stage___block_587_vnum2 = 0;
_t___block_592_cmp_yx = 0;
_t___block_592_cmp_zx = 0;
_t___block_592_cmp_zy = 0;
_t___block_592_x_sel = 0;
_t___block_592_y_sel = 0;
_t___block_592_z_sel = 0;
_t___stage___block_608_tex = 0;
_t___stage___block_608_vnum0 = 0;
_t___stage___block_608_vnum1 = 0;
_t___stage___block_608_vnum2 = 0;
_t___block_613_cmp_yx = 0;
_t___block_613_cmp_zx = 0;
_t___block_613_cmp_zy = 0;
_t___block_613_x_sel = 0;
_t___block_613_y_sel = 0;
_t___block_613_z_sel = 0;
_t___stage___block_629_tex = 0;
_t___stage___block_629_vnum0 = 0;
_t___stage___block_629_vnum1 = 0;
_t___stage___block_629_vnum2 = 0;
_t___block_634_cmp_yx = 0;
_t___block_634_cmp_zx = 0;
_t___block_634_cmp_zy = 0;
_t___block_634_x_sel = 0;
_t___block_634_y_sel = 0;
_t___block_634_z_sel = 0;
_t___stage___block_650_tex = 0;
_t___stage___block_650_vnum0 = 0;
_t___stage___block_650_vnum1 = 0;
_t___stage___block_650_vnum2 = 0;
_t___block_655_cmp_yx = 0;
_t___block_655_cmp_zx = 0;
_t___block_655_cmp_zy = 0;
_t___block_655_x_sel = 0;
_t___block_655_y_sel = 0;
_t___block_655_z_sel = 0;
_t___stage___block_671_tex = 0;
_t___stage___block_671_vnum0 = 0;
_t___stage___block_671_vnum1 = 0;
_t___stage___block_671_vnum2 = 0;
_t___block_676_cmp_yx = 0;
_t___block_676_cmp_zx = 0;
_t___block_676_cmp_zy = 0;
_t___block_676_x_sel = 0;
_t___block_676_y_sel = 0;
_t___block_676_z_sel = 0;
_t___stage___block_692_tex = 0;
_t___stage___block_692_vnum0 = 0;
_t___stage___block_692_vnum1 = 0;
_t___stage___block_692_vnum2 = 0;
_t___block_697_cmp_yx = 0;
_t___block_697_cmp_zx = 0;
_t___block_697_cmp_zy = 0;
_t___block_697_x_sel = 0;
_t___block_697_y_sel = 0;
_t___block_697_z_sel = 0;
_t___stage___block_713_tex = 0;
_t___stage___block_713_vnum0 = 0;
_t___stage___block_713_vnum1 = 0;
_t___stage___block_713_vnum2 = 0;
_t___block_718_cmp_yx = 0;
_t___block_718_cmp_zx = 0;
_t___block_718_cmp_zy = 0;
_t___block_718_x_sel = 0;
_t___block_718_y_sel = 0;
_t___block_718_z_sel = 0;
_t___stage___block_734_tex = 0;
_t___stage___block_734_vnum0 = 0;
_t___stage___block_734_vnum1 = 0;
_t___stage___block_734_vnum2 = 0;
_t___block_739_cmp_yx = 0;
_t___block_739_cmp_zx = 0;
_t___block_739_cmp_zy = 0;
_t___block_739_x_sel = 0;
_t___block_739_y_sel = 0;
_t___block_739_z_sel = 0;
_t___stage___block_755_tex = 0;
_t___stage___block_755_vnum0 = 0;
_t___stage___block_755_vnum1 = 0;
_t___stage___block_755_vnum2 = 0;
_t___block_760_cmp_yx = 0;
_t___block_760_cmp_zx = 0;
_t___block_760_cmp_zy = 0;
_t___block_760_x_sel = 0;
_t___block_760_y_sel = 0;
_t___block_760_z_sel = 0;
_t___stage___block_776_tex = 0;
_t___stage___block_776_vnum0 = 0;
_t___stage___block_776_vnum1 = 0;
_t___stage___block_776_vnum2 = 0;
_t___block_781_cmp_yx = 0;
_t___block_781_cmp_zx = 0;
_t___block_781_cmp_zy = 0;
_t___block_781_x_sel = 0;
_t___block_781_y_sel = 0;
_t___block_781_z_sel = 0;
_t___stage___block_797_tex = 0;
_t___stage___block_797_vnum0 = 0;
_t___stage___block_797_vnum1 = 0;
_t___stage___block_797_vnum2 = 0;
_t___block_802_cmp_yx = 0;
_t___block_802_cmp_zx = 0;
_t___block_802_cmp_zy = 0;
_t___block_802_x_sel = 0;
_t___block_802_y_sel = 0;
_t___block_802_z_sel = 0;
_t___stage___block_818_tex = 0;
_t___stage___block_818_vnum0 = 0;
_t___stage___block_818_vnum1 = 0;
_t___stage___block_818_vnum2 = 0;
_t___block_823_cmp_yx = 0;
_t___block_823_cmp_zx = 0;
_t___block_823_cmp_zy = 0;
_t___block_823_x_sel = 0;
_t___block_823_y_sel = 0;
_t___block_823_z_sel = 0;
_t___stage___block_839_tex = 0;
_t___stage___block_839_vnum0 = 0;
_t___stage___block_839_vnum1 = 0;
_t___stage___block_839_vnum2 = 0;
_t___block_844_cmp_yx = 0;
_t___block_844_cmp_zx = 0;
_t___block_844_cmp_zy = 0;
_t___block_844_x_sel = 0;
_t___block_844_y_sel = 0;
_t___block_844_z_sel = 0;
_t___stage___block_860_tex = 0;
_t___stage___block_860_vnum0 = 0;
_t___stage___block_860_vnum1 = 0;
_t___stage___block_860_vnum2 = 0;
_t___block_865_cmp_yx = 0;
_t___block_865_cmp_zx = 0;
_t___block_865_cmp_zy = 0;
_t___block_865_x_sel = 0;
_t___block_865_y_sel = 0;
_t___block_865_z_sel = 0;
_t___stage___block_881_tex = 0;
_t___stage___block_881_vnum0 = 0;
_t___stage___block_881_vnum1 = 0;
_t___stage___block_881_vnum2 = 0;
_t___block_886_cmp_yx = 0;
_t___block_886_cmp_zx = 0;
_t___block_886_cmp_zy = 0;
_t___block_886_x_sel = 0;
_t___block_886_y_sel = 0;
_t___block_886_z_sel = 0;
_t___stage___block_902_tex = 0;
_t___stage___block_902_vnum0 = 0;
_t___stage___block_902_vnum1 = 0;
_t___stage___block_902_vnum2 = 0;
_t___block_907_cmp_yx = 0;
_t___block_907_cmp_zx = 0;
_t___block_907_cmp_zy = 0;
_t___block_907_x_sel = 0;
_t___block_907_y_sel = 0;
_t___block_907_z_sel = 0;
_t___stage___block_923_tex = 0;
_t___stage___block_923_vnum0 = 0;
_t___stage___block_923_vnum1 = 0;
_t___stage___block_923_vnum2 = 0;
_t___block_928_cmp_yx = 0;
_t___block_928_cmp_zx = 0;
_t___block_928_cmp_zy = 0;
_t___block_928_x_sel = 0;
_t___block_928_y_sel = 0;
_t___block_928_z_sel = 0;
_t___stage___block_944_tex = 0;
_t___stage___block_944_vnum0 = 0;
_t___stage___block_944_vnum1 = 0;
_t___stage___block_944_vnum2 = 0;
_t___block_949_cmp_yx = 0;
_t___block_949_cmp_zx = 0;
_t___block_949_cmp_zy = 0;
_t___block_949_x_sel = 0;
_t___block_949_y_sel = 0;
_t___block_949_z_sel = 0;
_t___stage___block_965_tex = 0;
_t___stage___block_965_vnum0 = 0;
_t___stage___block_965_vnum1 = 0;
_t___stage___block_965_vnum2 = 0;
_t___block_970_cmp_yx = 0;
_t___block_970_cmp_zx = 0;
_t___block_970_cmp_zy = 0;
_t___block_970_x_sel = 0;
_t___block_970_y_sel = 0;
_t___block_970_z_sel = 0;
_t___stage___block_986_tex = 0;
_t___stage___block_986_vnum0 = 0;
_t___stage___block_986_vnum1 = 0;
_t___stage___block_986_vnum2 = 0;
_t___block_991_cmp_yx = 0;
_t___block_991_cmp_zx = 0;
_t___block_991_cmp_zy = 0;
_t___block_991_x_sel = 0;
_t___block_991_y_sel = 0;
_t___block_991_z_sel = 0;
_t___stage___block_1007_tex = 0;
_t___stage___block_1007_vnum0 = 0;
_t___stage___block_1007_vnum1 = 0;
_t___stage___block_1007_vnum2 = 0;
_t___block_1012_cmp_yx = 0;
_t___block_1012_cmp_zx = 0;
_t___block_1012_cmp_zy = 0;
_t___block_1012_x_sel = 0;
_t___block_1012_y_sel = 0;
_t___block_1012_z_sel = 0;
_t___stage___block_1028_tex = 0;
_t___stage___block_1028_vnum0 = 0;
_t___stage___block_1028_vnum1 = 0;
_t___stage___block_1028_vnum2 = 0;
_t___block_1033_cmp_yx = 0;
_t___block_1033_cmp_zx = 0;
_t___block_1033_cmp_zy = 0;
_t___block_1033_x_sel = 0;
_t___block_1033_y_sel = 0;
_t___block_1033_z_sel = 0;
_t___stage___block_1049_tex = 0;
_t___stage___block_1049_vnum0 = 0;
_t___stage___block_1049_vnum1 = 0;
_t___stage___block_1049_vnum2 = 0;
_t___block_1054_cmp_yx = 0;
_t___block_1054_cmp_zx = 0;
_t___block_1054_cmp_zy = 0;
_t___block_1054_x_sel = 0;
_t___block_1054_y_sel = 0;
_t___block_1054_z_sel = 0;
_t___stage___block_1070_tex = 0;
_t___stage___block_1070_vnum0 = 0;
_t___stage___block_1070_vnum1 = 0;
_t___stage___block_1070_vnum2 = 0;
_t___block_1075_cmp_yx = 0;
_t___block_1075_cmp_zx = 0;
_t___block_1075_cmp_zy = 0;
_t___block_1075_x_sel = 0;
_t___block_1075_y_sel = 0;
_t___block_1075_z_sel = 0;
_t___stage___block_1091_tex = 0;
_t___stage___block_1091_vnum0 = 0;
_t___stage___block_1091_vnum1 = 0;
_t___stage___block_1091_vnum2 = 0;
_t___block_1096_cmp_yx = 0;
_t___block_1096_cmp_zx = 0;
_t___block_1096_cmp_zy = 0;
_t___block_1096_x_sel = 0;
_t___block_1096_y_sel = 0;
_t___block_1096_z_sel = 0;
_t___stage___block_1112_tex = 0;
_t___stage___block_1112_vnum0 = 0;
_t___stage___block_1112_vnum1 = 0;
_t___stage___block_1112_vnum2 = 0;
_t___block_1117_cmp_yx = 0;
_t___block_1117_cmp_zx = 0;
_t___block_1117_cmp_zy = 0;
_t___block_1117_x_sel = 0;
_t___block_1117_y_sel = 0;
_t___block_1117_z_sel = 0;
_t___stage___block_1133_tex = 0;
_t___stage___block_1133_vnum0 = 0;
_t___stage___block_1133_vnum1 = 0;
_t___stage___block_1133_vnum2 = 0;
_t___block_1138_cmp_yx = 0;
_t___block_1138_cmp_zx = 0;
_t___block_1138_cmp_zy = 0;
_t___block_1138_x_sel = 0;
_t___block_1138_y_sel = 0;
_t___block_1138_z_sel = 0;
_t___stage___block_1154_tex = 0;
_t___stage___block_1154_vnum0 = 0;
_t___stage___block_1154_vnum1 = 0;
_t___stage___block_1154_vnum2 = 0;
_t___block_1159_cmp_yx = 0;
_t___block_1159_cmp_zx = 0;
_t___block_1159_cmp_zy = 0;
_t___block_1159_x_sel = 0;
_t___block_1159_y_sel = 0;
_t___block_1159_z_sel = 0;
_t___stage___block_1175_tex = 0;
_t___stage___block_1175_vnum0 = 0;
_t___stage___block_1175_vnum1 = 0;
_t___stage___block_1175_vnum2 = 0;
_t___block_1180_cmp_yx = 0;
_t___block_1180_cmp_zx = 0;
_t___block_1180_cmp_zy = 0;
_t___block_1180_x_sel = 0;
_t___block_1180_y_sel = 0;
_t___block_1180_z_sel = 0;
_t___stage___block_1196_tex = 0;
_t___stage___block_1196_vnum0 = 0;
_t___stage___block_1196_vnum1 = 0;
_t___stage___block_1196_vnum2 = 0;
_t___block_1201_cmp_yx = 0;
_t___block_1201_cmp_zx = 0;
_t___block_1201_cmp_zy = 0;
_t___block_1201_x_sel = 0;
_t___block_1201_y_sel = 0;
_t___block_1201_z_sel = 0;
_t___stage___block_1217_tex = 0;
_t___stage___block_1217_vnum0 = 0;
_t___stage___block_1217_vnum1 = 0;
_t___stage___block_1217_vnum2 = 0;
_t___block_1222_cmp_yx = 0;
_t___block_1222_cmp_zx = 0;
_t___block_1222_cmp_zy = 0;
_t___block_1222_x_sel = 0;
_t___block_1222_y_sel = 0;
_t___block_1222_z_sel = 0;
_t___stage___block_1238_tex = 0;
_t___stage___block_1238_vnum0 = 0;
_t___stage___block_1238_vnum1 = 0;
_t___stage___block_1238_vnum2 = 0;
_t___block_1243_cmp_yx = 0;
_t___block_1243_cmp_zx = 0;
_t___block_1243_cmp_zy = 0;
_t___block_1243_x_sel = 0;
_t___block_1243_y_sel = 0;
_t___block_1243_z_sel = 0;
_t___stage___block_1259_tex = 0;
_t___stage___block_1259_vnum0 = 0;
_t___stage___block_1259_vnum1 = 0;
_t___stage___block_1259_vnum2 = 0;
_t___block_1264_cmp_yx = 0;
_t___block_1264_cmp_zx = 0;
_t___block_1264_cmp_zy = 0;
_t___block_1264_x_sel = 0;
_t___block_1264_y_sel = 0;
_t___block_1264_z_sel = 0;
_t___stage___block_1280_tex = 0;
_t___stage___block_1280_vnum0 = 0;
_t___stage___block_1280_vnum1 = 0;
_t___stage___block_1280_vnum2 = 0;
_t___block_1285_cmp_yx = 0;
_t___block_1285_cmp_zx = 0;
_t___block_1285_cmp_zy = 0;
_t___block_1285_x_sel = 0;
_t___block_1285_y_sel = 0;
_t___block_1285_z_sel = 0;
_t___stage___block_1301_tex = 0;
_t___stage___block_1301_vnum0 = 0;
_t___stage___block_1301_vnum1 = 0;
_t___stage___block_1301_vnum2 = 0;
_t___block_1306_cmp_yx = 0;
_t___block_1306_cmp_zx = 0;
_t___block_1306_cmp_zy = 0;
_t___block_1306_x_sel = 0;
_t___block_1306_y_sel = 0;
_t___block_1306_z_sel = 0;
_t___stage___block_1322_tex = 0;
_t___stage___block_1322_vnum0 = 0;
_t___stage___block_1322_vnum1 = 0;
_t___stage___block_1322_vnum2 = 0;
_t___block_1327_cmp_yx = 0;
_t___block_1327_cmp_zx = 0;
_t___block_1327_cmp_zy = 0;
_t___block_1327_x_sel = 0;
_t___block_1327_y_sel = 0;
_t___block_1327_z_sel = 0;
_t___stage___block_1343_tex = 0;
_t___stage___block_1343_vnum0 = 0;
_t___stage___block_1343_vnum1 = 0;
_t___stage___block_1343_vnum2 = 0;
_t___block_1348_cmp_yx = 0;
_t___block_1348_cmp_zx = 0;
_t___block_1348_cmp_zy = 0;
_t___block_1348_x_sel = 0;
_t___block_1348_y_sel = 0;
_t___block_1348_z_sel = 0;
_t___stage___block_1364_tex = 0;
_t___stage___block_1364_vnum0 = 0;
_t___stage___block_1364_vnum1 = 0;
_t___stage___block_1364_vnum2 = 0;
_t___block_1369_cmp_yx = 0;
_t___block_1369_cmp_zx = 0;
_t___block_1369_cmp_zy = 0;
_t___block_1369_x_sel = 0;
_t___block_1369_y_sel = 0;
_t___block_1369_z_sel = 0;
_t___stage___block_1385_tex = 0;
_t___stage___block_1385_vnum0 = 0;
_t___stage___block_1385_vnum1 = 0;
_t___stage___block_1385_vnum2 = 0;
_t___block_1390_cmp_yx = 0;
_t___block_1390_cmp_zx = 0;
_t___block_1390_cmp_zy = 0;
_t___block_1390_x_sel = 0;
_t___block_1390_y_sel = 0;
_t___block_1390_z_sel = 0;
_t___stage___block_1406_tex = 0;
_t___stage___block_1406_vnum0 = 0;
_t___stage___block_1406_vnum1 = 0;
_t___stage___block_1406_vnum2 = 0;
_t___block_1411_cmp_yx = 0;
_t___block_1411_cmp_zx = 0;
_t___block_1411_cmp_zy = 0;
_t___block_1411_x_sel = 0;
_t___block_1411_y_sel = 0;
_t___block_1411_z_sel = 0;
_t___stage___block_1427_tex = 0;
_t___stage___block_1427_vnum0 = 0;
_t___stage___block_1427_vnum1 = 0;
_t___stage___block_1427_vnum2 = 0;
_t___block_1432_cmp_yx = 0;
_t___block_1432_cmp_zx = 0;
_t___block_1432_cmp_zy = 0;
_t___block_1432_x_sel = 0;
_t___block_1432_y_sel = 0;
_t___block_1432_z_sel = 0;
_t___stage___block_1448_tex = 0;
_t___stage___block_1448_vnum0 = 0;
_t___stage___block_1448_vnum1 = 0;
_t___stage___block_1448_vnum2 = 0;
_t___block_1453_cmp_yx = 0;
_t___block_1453_cmp_zx = 0;
_t___block_1453_cmp_zy = 0;
_t___block_1453_x_sel = 0;
_t___block_1453_y_sel = 0;
_t___block_1453_z_sel = 0;
_t___stage___block_1469_tex = 0;
_t___stage___block_1469_vnum0 = 0;
_t___stage___block_1469_vnum1 = 0;
_t___stage___block_1469_vnum2 = 0;
_t___block_1474_cmp_yx = 0;
_t___block_1474_cmp_zx = 0;
_t___block_1474_cmp_zy = 0;
_t___block_1474_x_sel = 0;
_t___block_1474_y_sel = 0;
_t___block_1474_z_sel = 0;
_t___stage___block_1490_tex = 0;
_t___stage___block_1490_vnum0 = 0;
_t___stage___block_1490_vnum1 = 0;
_t___stage___block_1490_vnum2 = 0;
_t___block_1495_cmp_yx = 0;
_t___block_1495_cmp_zx = 0;
_t___block_1495_cmp_zy = 0;
_t___block_1495_x_sel = 0;
_t___block_1495_y_sel = 0;
_t___block_1495_z_sel = 0;
_t___stage___block_1511_tex = 0;
_t___stage___block_1511_vnum0 = 0;
_t___stage___block_1511_vnum1 = 0;
_t___stage___block_1511_vnum2 = 0;
_t___block_1516_cmp_yx = 0;
_t___block_1516_cmp_zx = 0;
_t___block_1516_cmp_zy = 0;
_t___block_1516_x_sel = 0;
_t___block_1516_y_sel = 0;
_t___block_1516_z_sel = 0;
_t___stage___block_1532_tex = 0;
_t___stage___block_1532_vnum0 = 0;
_t___stage___block_1532_vnum1 = 0;
_t___stage___block_1532_vnum2 = 0;
_t___block_1537_cmp_yx = 0;
_t___block_1537_cmp_zx = 0;
_t___block_1537_cmp_zy = 0;
_t___block_1537_x_sel = 0;
_t___block_1537_y_sel = 0;
_t___block_1537_z_sel = 0;
_t___stage___block_1553_tex = 0;
_t___stage___block_1553_vnum0 = 0;
_t___stage___block_1553_vnum1 = 0;
_t___stage___block_1553_vnum2 = 0;
_t___block_1558_cmp_yx = 0;
_t___block_1558_cmp_zx = 0;
_t___block_1558_cmp_zy = 0;
_t___block_1558_x_sel = 0;
_t___block_1558_y_sel = 0;
_t___block_1558_z_sel = 0;
_t___stage___block_1574_tex = 0;
_t___stage___block_1574_vnum0 = 0;
_t___stage___block_1574_vnum1 = 0;
_t___stage___block_1574_vnum2 = 0;
_t___block_1579_cmp_yx = 0;
_t___block_1579_cmp_zx = 0;
_t___block_1579_cmp_zy = 0;
_t___block_1579_x_sel = 0;
_t___block_1579_y_sel = 0;
_t___block_1579_z_sel = 0;
_t___stage___block_1595_tex = 0;
_t___stage___block_1595_vnum0 = 0;
_t___stage___block_1595_vnum1 = 0;
_t___stage___block_1595_vnum2 = 0;
_t___block_1600_cmp_yx = 0;
_t___block_1600_cmp_zx = 0;
_t___block_1600_cmp_zy = 0;
_t___block_1600_x_sel = 0;
_t___block_1600_y_sel = 0;
_t___block_1600_z_sel = 0;
_t___stage___block_1616_tex = 0;
_t___stage___block_1616_vnum0 = 0;
_t___stage___block_1616_vnum1 = 0;
_t___stage___block_1616_vnum2 = 0;
_t___block_1621_cmp_yx = 0;
_t___block_1621_cmp_zx = 0;
_t___block_1621_cmp_zy = 0;
_t___block_1621_x_sel = 0;
_t___block_1621_y_sel = 0;
_t___block_1621_z_sel = 0;
_t___stage___block_1637_tex = 0;
_t___stage___block_1637_vnum0 = 0;
_t___stage___block_1637_vnum1 = 0;
_t___stage___block_1637_vnum2 = 0;
_t___block_1642_cmp_yx = 0;
_t___block_1642_cmp_zx = 0;
_t___block_1642_cmp_zy = 0;
_t___block_1642_x_sel = 0;
_t___block_1642_y_sel = 0;
_t___block_1642_z_sel = 0;
_t___stage___block_1658_tex = 0;
_t___stage___block_1658_vnum0 = 0;
_t___stage___block_1658_vnum1 = 0;
_t___stage___block_1658_vnum2 = 0;
_t___block_1663_cmp_yx = 0;
_t___block_1663_cmp_zx = 0;
_t___block_1663_cmp_zy = 0;
_t___block_1663_x_sel = 0;
_t___block_1663_y_sel = 0;
_t___block_1663_z_sel = 0;
_t___stage___block_1679_tex = 0;
_t___stage___block_1679_vnum0 = 0;
_t___stage___block_1679_vnum1 = 0;
_t___stage___block_1679_vnum2 = 0;
_t___block_1684_cmp_yx = 0;
_t___block_1684_cmp_zx = 0;
_t___block_1684_cmp_zy = 0;
_t___block_1684_x_sel = 0;
_t___block_1684_y_sel = 0;
_t___block_1684_z_sel = 0;
_t___stage___block_1700_tex = 0;
_t___stage___block_1700_vnum0 = 0;
_t___stage___block_1700_vnum1 = 0;
_t___stage___block_1700_vnum2 = 0;
_t___block_1705_cmp_yx = 0;
_t___block_1705_cmp_zx = 0;
_t___block_1705_cmp_zy = 0;
_t___block_1705_x_sel = 0;
_t___block_1705_y_sel = 0;
_t___block_1705_z_sel = 0;
_t___stage___block_1721_tex = 0;
_t___stage___block_1721_vnum0 = 0;
_t___stage___block_1721_vnum1 = 0;
_t___stage___block_1721_vnum2 = 0;
_t___block_1726_cmp_yx = 0;
_t___block_1726_cmp_zx = 0;
_t___block_1726_cmp_zy = 0;
_t___block_1726_x_sel = 0;
_t___block_1726_y_sel = 0;
_t___block_1726_z_sel = 0;
_t___stage___block_1742_tex = 0;
_t___stage___block_1742_vnum0 = 0;
_t___stage___block_1742_vnum1 = 0;
_t___stage___block_1742_vnum2 = 0;
_t___block_1747_cmp_yx = 0;
_t___block_1747_cmp_zx = 0;
_t___block_1747_cmp_zy = 0;
_t___block_1747_x_sel = 0;
_t___block_1747_y_sel = 0;
_t___block_1747_z_sel = 0;
_t___stage___block_1763_tex = 0;
_t___stage___block_1763_vnum0 = 0;
_t___stage___block_1763_vnum1 = 0;
_t___stage___block_1763_vnum2 = 0;
_t___block_1768_cmp_yx = 0;
_t___block_1768_cmp_zx = 0;
_t___block_1768_cmp_zy = 0;
_t___block_1768_x_sel = 0;
_t___block_1768_y_sel = 0;
_t___block_1768_z_sel = 0;
_t___stage___block_1784_tex = 0;
_t___stage___block_1784_vnum0 = 0;
_t___stage___block_1784_vnum1 = 0;
_t___stage___block_1784_vnum2 = 0;
_t___block_1789_cmp_yx = 0;
_t___block_1789_cmp_zx = 0;
_t___block_1789_cmp_zy = 0;
_t___block_1789_x_sel = 0;
_t___block_1789_y_sel = 0;
_t___block_1789_z_sel = 0;
_t___stage___block_1805_tex = 0;
_t___stage___block_1805_vnum0 = 0;
_t___stage___block_1805_vnum1 = 0;
_t___stage___block_1805_vnum2 = 0;
_t___block_1810_cmp_yx = 0;
_t___block_1810_cmp_zx = 0;
_t___block_1810_cmp_zy = 0;
_t___block_1810_x_sel = 0;
_t___block_1810_y_sel = 0;
_t___block_1810_z_sel = 0;
_t___stage___block_1826_tex = 0;
_t___stage___block_1826_vnum0 = 0;
_t___stage___block_1826_vnum1 = 0;
_t___stage___block_1826_vnum2 = 0;
_t___block_1831_cmp_yx = 0;
_t___block_1831_cmp_zx = 0;
_t___block_1831_cmp_zy = 0;
_t___block_1831_x_sel = 0;
_t___block_1831_y_sel = 0;
_t___block_1831_z_sel = 0;
_t___stage___block_1847_tex = 0;
_t___stage___block_1847_vnum0 = 0;
_t___stage___block_1847_vnum1 = 0;
_t___stage___block_1847_vnum2 = 0;
_t___block_1852_cmp_yx = 0;
_t___block_1852_cmp_zx = 0;
_t___block_1852_cmp_zy = 0;
_t___block_1852_x_sel = 0;
_t___block_1852_y_sel = 0;
_t___block_1852_z_sel = 0;
_t___stage___block_1868_tex = 0;
_t___stage___block_1868_vnum0 = 0;
_t___stage___block_1868_vnum1 = 0;
_t___stage___block_1868_vnum2 = 0;
_t___block_1873_cmp_yx = 0;
_t___block_1873_cmp_zx = 0;
_t___block_1873_cmp_zy = 0;
_t___block_1873_x_sel = 0;
_t___block_1873_y_sel = 0;
_t___block_1873_z_sel = 0;
_t___stage___block_1889_tex = 0;
_t___stage___block_1889_vnum0 = 0;
_t___stage___block_1889_vnum1 = 0;
_t___stage___block_1889_vnum2 = 0;
_t___block_1894_cmp_yx = 0;
_t___block_1894_cmp_zx = 0;
_t___block_1894_cmp_zy = 0;
_t___block_1894_x_sel = 0;
_t___block_1894_y_sel = 0;
_t___block_1894_z_sel = 0;
_t___stage___block_1910_tex = 0;
_t___stage___block_1910_vnum0 = 0;
_t___stage___block_1910_vnum1 = 0;
_t___stage___block_1910_vnum2 = 0;
_t___block_1915_cmp_yx = 0;
_t___block_1915_cmp_zx = 0;
_t___block_1915_cmp_zy = 0;
_t___block_1915_x_sel = 0;
_t___block_1915_y_sel = 0;
_t___block_1915_z_sel = 0;
_t___stage___block_1931_tex = 0;
_t___stage___block_1931_vnum0 = 0;
_t___stage___block_1931_vnum1 = 0;
_t___stage___block_1931_vnum2 = 0;
_t___block_1936_cmp_yx = 0;
_t___block_1936_cmp_zx = 0;
_t___block_1936_cmp_zy = 0;
_t___block_1936_x_sel = 0;
_t___block_1936_y_sel = 0;
_t___block_1936_z_sel = 0;
_t___stage___block_1952_tex = 0;
_t___stage___block_1952_vnum0 = 0;
_t___stage___block_1952_vnum1 = 0;
_t___stage___block_1952_vnum2 = 0;
_t___block_1957_cmp_yx = 0;
_t___block_1957_cmp_zx = 0;
_t___block_1957_cmp_zy = 0;
_t___block_1957_x_sel = 0;
_t___block_1957_y_sel = 0;
_t___block_1957_z_sel = 0;
_t___stage___block_1973_tex = 0;
_t___stage___block_1973_vnum0 = 0;
_t___stage___block_1973_vnum1 = 0;
_t___stage___block_1973_vnum2 = 0;
_t___block_1978_cmp_yx = 0;
_t___block_1978_cmp_zx = 0;
_t___block_1978_cmp_zy = 0;
_t___block_1978_x_sel = 0;
_t___block_1978_y_sel = 0;
_t___block_1978_z_sel = 0;
_t___stage___block_1994_tex = 0;
_t___stage___block_1994_vnum0 = 0;
_t___stage___block_1994_vnum1 = 0;
_t___stage___block_1994_vnum2 = 0;
_t___block_1999_cmp_yx = 0;
_t___block_1999_cmp_zx = 0;
_t___block_1999_cmp_zy = 0;
_t___block_1999_x_sel = 0;
_t___block_1999_y_sel = 0;
_t___block_1999_z_sel = 0;
_t___stage___block_2015_tex = 0;
_t___stage___block_2015_vnum0 = 0;
_t___stage___block_2015_vnum1 = 0;
_t___stage___block_2015_vnum2 = 0;
_t___block_2020_cmp_yx = 0;
_t___block_2020_cmp_zx = 0;
_t___block_2020_cmp_zy = 0;
_t___block_2020_x_sel = 0;
_t___block_2020_y_sel = 0;
_t___block_2020_z_sel = 0;
_t___stage___block_2036_tex = 0;
_t___stage___block_2036_vnum0 = 0;
_t___stage___block_2036_vnum1 = 0;
_t___stage___block_2036_vnum2 = 0;
_t___block_2041_cmp_yx = 0;
_t___block_2041_cmp_zx = 0;
_t___block_2041_cmp_zy = 0;
_t___block_2041_x_sel = 0;
_t___block_2041_y_sel = 0;
_t___block_2041_z_sel = 0;
_t___stage___block_2057_tex = 0;
_t___stage___block_2057_vnum0 = 0;
_t___stage___block_2057_vnum1 = 0;
_t___stage___block_2057_vnum2 = 0;
_t___block_2062_cmp_yx = 0;
_t___block_2062_cmp_zx = 0;
_t___block_2062_cmp_zy = 0;
_t___block_2062_x_sel = 0;
_t___block_2062_y_sel = 0;
_t___block_2062_z_sel = 0;
_t___stage___block_2078_tex = 0;
_t___stage___block_2078_vnum0 = 0;
_t___stage___block_2078_vnum1 = 0;
_t___stage___block_2078_vnum2 = 0;
_t___block_2083_cmp_yx = 0;
_t___block_2083_cmp_zx = 0;
_t___block_2083_cmp_zy = 0;
_t___block_2083_x_sel = 0;
_t___block_2083_y_sel = 0;
_t___block_2083_z_sel = 0;
_t___stage___block_2099_tex = 0;
_t___stage___block_2099_vnum0 = 0;
_t___stage___block_2099_vnum1 = 0;
_t___stage___block_2099_vnum2 = 0;
_t___block_2104_cmp_yx = 0;
_t___block_2104_cmp_zx = 0;
_t___block_2104_cmp_zy = 0;
_t___block_2104_x_sel = 0;
_t___block_2104_y_sel = 0;
_t___block_2104_z_sel = 0;
_t___stage___block_2120_tex = 0;
_t___stage___block_2120_vnum0 = 0;
_t___stage___block_2120_vnum1 = 0;
_t___stage___block_2120_vnum2 = 0;
_t___block_2125_cmp_yx = 0;
_t___block_2125_cmp_zx = 0;
_t___block_2125_cmp_zy = 0;
_t___block_2125_x_sel = 0;
_t___block_2125_y_sel = 0;
_t___block_2125_z_sel = 0;
_t___stage___block_2141_tex = 0;
_t___stage___block_2141_vnum0 = 0;
_t___stage___block_2141_vnum1 = 0;
_t___stage___block_2141_vnum2 = 0;
_t___block_2146_cmp_yx = 0;
_t___block_2146_cmp_zx = 0;
_t___block_2146_cmp_zy = 0;
_t___block_2146_x_sel = 0;
_t___block_2146_y_sel = 0;
_t___block_2146_z_sel = 0;
_t___stage___block_2162_tex = 0;
_t___stage___block_2162_vnum0 = 0;
_t___stage___block_2162_vnum1 = 0;
_t___stage___block_2162_vnum2 = 0;
_t___block_2167_cmp_yx = 0;
_t___block_2167_cmp_zx = 0;
_t___block_2167_cmp_zy = 0;
_t___block_2167_x_sel = 0;
_t___block_2167_y_sel = 0;
_t___block_2167_z_sel = 0;
_t___stage___block_2183_tex = 0;
_t___stage___block_2183_vnum0 = 0;
_t___stage___block_2183_vnum1 = 0;
_t___stage___block_2183_vnum2 = 0;
_t___block_2188_cmp_yx = 0;
_t___block_2188_cmp_zx = 0;
_t___block_2188_cmp_zy = 0;
_t___block_2188_x_sel = 0;
_t___block_2188_y_sel = 0;
_t___block_2188_z_sel = 0;
_t___stage___block_2204_tex = 0;
_t___stage___block_2204_vnum0 = 0;
_t___stage___block_2204_vnum1 = 0;
_t___stage___block_2204_vnum2 = 0;
_t___block_2209_cmp_yx = 0;
_t___block_2209_cmp_zx = 0;
_t___block_2209_cmp_zy = 0;
_t___block_2209_x_sel = 0;
_t___block_2209_y_sel = 0;
_t___block_2209_z_sel = 0;
_t___stage___block_2225_tex = 0;
_t___stage___block_2225_vnum0 = 0;
_t___stage___block_2225_vnum1 = 0;
_t___stage___block_2225_vnum2 = 0;
_t___block_2230_cmp_yx = 0;
_t___block_2230_cmp_zx = 0;
_t___block_2230_cmp_zy = 0;
_t___block_2230_x_sel = 0;
_t___block_2230_y_sel = 0;
_t___block_2230_z_sel = 0;
_t___stage___block_2246_tex = 0;
_t___stage___block_2246_vnum0 = 0;
_t___stage___block_2246_vnum1 = 0;
_t___stage___block_2246_vnum2 = 0;
_t___block_2251_cmp_yx = 0;
_t___block_2251_cmp_zx = 0;
_t___block_2251_cmp_zy = 0;
_t___block_2251_x_sel = 0;
_t___block_2251_y_sel = 0;
_t___block_2251_z_sel = 0;
_t___stage___block_2267_tex = 0;
_t___stage___block_2267_vnum0 = 0;
_t___stage___block_2267_vnum1 = 0;
_t___stage___block_2267_vnum2 = 0;
_t___block_2272_cmp_yx = 0;
_t___block_2272_cmp_zx = 0;
_t___block_2272_cmp_zy = 0;
_t___block_2272_x_sel = 0;
_t___block_2272_y_sel = 0;
_t___block_2272_z_sel = 0;
_t___stage___block_2288_tex = 0;
_t___stage___block_2288_vnum0 = 0;
_t___stage___block_2288_vnum1 = 0;
_t___stage___block_2288_vnum2 = 0;
_t___block_2293_cmp_yx = 0;
_t___block_2293_cmp_zx = 0;
_t___block_2293_cmp_zy = 0;
_t___block_2293_x_sel = 0;
_t___block_2293_y_sel = 0;
_t___block_2293_z_sel = 0;
_t___stage___block_2309_tex = 0;
_t___stage___block_2309_vnum0 = 0;
_t___stage___block_2309_vnum1 = 0;
_t___stage___block_2309_vnum2 = 0;
_t___block_2314_cmp_yx = 0;
_t___block_2314_cmp_zx = 0;
_t___block_2314_cmp_zy = 0;
_t___block_2314_x_sel = 0;
_t___block_2314_y_sel = 0;
_t___block_2314_z_sel = 0;
_t___stage___block_2330_tex = 0;
_t___stage___block_2330_vnum0 = 0;
_t___stage___block_2330_vnum1 = 0;
_t___stage___block_2330_vnum2 = 0;
_t___block_2335_cmp_yx = 0;
_t___block_2335_cmp_zx = 0;
_t___block_2335_cmp_zy = 0;
_t___block_2335_x_sel = 0;
_t___block_2335_y_sel = 0;
_t___block_2335_z_sel = 0;
_t___stage___block_2351_tex = 0;
_t___stage___block_2351_vnum0 = 0;
_t___stage___block_2351_vnum1 = 0;
_t___stage___block_2351_vnum2 = 0;
_t___block_2356_cmp_yx = 0;
_t___block_2356_cmp_zx = 0;
_t___block_2356_cmp_zy = 0;
_t___block_2356_x_sel = 0;
_t___block_2356_y_sel = 0;
_t___block_2356_z_sel = 0;
_t___stage___block_2372_tex = 0;
_t___stage___block_2372_vnum0 = 0;
_t___stage___block_2372_vnum1 = 0;
_t___stage___block_2372_vnum2 = 0;
_t___block_2377_cmp_yx = 0;
_t___block_2377_cmp_zx = 0;
_t___block_2377_cmp_zy = 0;
_t___block_2377_x_sel = 0;
_t___block_2377_y_sel = 0;
_t___block_2377_z_sel = 0;
_t___stage___block_2393_tex = 0;
_t___stage___block_2393_vnum0 = 0;
_t___stage___block_2393_vnum1 = 0;
_t___stage___block_2393_vnum2 = 0;
_t___block_2398_cmp_yx = 0;
_t___block_2398_cmp_zx = 0;
_t___block_2398_cmp_zy = 0;
_t___block_2398_x_sel = 0;
_t___block_2398_y_sel = 0;
_t___block_2398_z_sel = 0;
_t___stage___block_2414_tex = 0;
_t___stage___block_2414_vnum0 = 0;
_t___stage___block_2414_vnum1 = 0;
_t___stage___block_2414_vnum2 = 0;
_t___block_2419_cmp_yx = 0;
_t___block_2419_cmp_zx = 0;
_t___block_2419_cmp_zy = 0;
_t___block_2419_x_sel = 0;
_t___block_2419_y_sel = 0;
_t___block_2419_z_sel = 0;
_t___stage___block_2435_tex = 0;
_t___stage___block_2435_vnum0 = 0;
_t___stage___block_2435_vnum1 = 0;
_t___stage___block_2435_vnum2 = 0;
_t___block_2440_cmp_yx = 0;
_t___block_2440_cmp_zx = 0;
_t___block_2440_cmp_zy = 0;
_t___block_2440_x_sel = 0;
_t___block_2440_y_sel = 0;
_t___block_2440_z_sel = 0;
_t___stage___block_2456_tex = 0;
_t___stage___block_2456_vnum0 = 0;
_t___stage___block_2456_vnum1 = 0;
_t___stage___block_2456_vnum2 = 0;
_t___block_2461_cmp_yx = 0;
_t___block_2461_cmp_zx = 0;
_t___block_2461_cmp_zy = 0;
_t___block_2461_x_sel = 0;
_t___block_2461_y_sel = 0;
_t___block_2461_z_sel = 0;
_t___stage___block_2477_tex = 0;
_t___stage___block_2477_vnum0 = 0;
_t___stage___block_2477_vnum1 = 0;
_t___stage___block_2477_vnum2 = 0;
_t___block_2482_cmp_yx = 0;
_t___block_2482_cmp_zx = 0;
_t___block_2482_cmp_zy = 0;
_t___block_2482_x_sel = 0;
_t___block_2482_y_sel = 0;
_t___block_2482_z_sel = 0;
_t___stage___block_2498_tex = 0;
_t___stage___block_2498_vnum0 = 0;
_t___stage___block_2498_vnum1 = 0;
_t___stage___block_2498_vnum2 = 0;
_t___block_2503_cmp_yx = 0;
_t___block_2503_cmp_zx = 0;
_t___block_2503_cmp_zy = 0;
_t___block_2503_x_sel = 0;
_t___block_2503_y_sel = 0;
_t___block_2503_z_sel = 0;
_t___stage___block_2519_tex = 0;
_t___stage___block_2519_vnum0 = 0;
_t___stage___block_2519_vnum1 = 0;
_t___stage___block_2519_vnum2 = 0;
_t___block_2524_cmp_yx = 0;
_t___block_2524_cmp_zx = 0;
_t___block_2524_cmp_zy = 0;
_t___block_2524_x_sel = 0;
_t___block_2524_y_sel = 0;
_t___block_2524_z_sel = 0;
_t___stage___block_2540_tex = 0;
_t___stage___block_2540_vnum0 = 0;
_t___stage___block_2540_vnum1 = 0;
_t___stage___block_2540_vnum2 = 0;
_t___block_2545_cmp_yx = 0;
_t___block_2545_cmp_zx = 0;
_t___block_2545_cmp_zy = 0;
_t___block_2545_x_sel = 0;
_t___block_2545_y_sel = 0;
_t___block_2545_z_sel = 0;
_t___stage___block_2561_tex = 0;
_t___stage___block_2561_vnum0 = 0;
_t___stage___block_2561_vnum1 = 0;
_t___stage___block_2561_vnum2 = 0;
_t___block_2566_cmp_yx = 0;
_t___block_2566_cmp_zx = 0;
_t___block_2566_cmp_zy = 0;
_t___block_2566_x_sel = 0;
_t___block_2566_y_sel = 0;
_t___block_2566_z_sel = 0;
_t___stage___block_2582_tex = 0;
_t___stage___block_2582_vnum0 = 0;
_t___stage___block_2582_vnum1 = 0;
_t___stage___block_2582_vnum2 = 0;
_t___block_2587_cmp_yx = 0;
_t___block_2587_cmp_zx = 0;
_t___block_2587_cmp_zy = 0;
_t___block_2587_x_sel = 0;
_t___block_2587_y_sel = 0;
_t___block_2587_z_sel = 0;
_t___stage___block_2603_tex = 0;
_t___stage___block_2603_vnum0 = 0;
_t___stage___block_2603_vnum1 = 0;
_t___stage___block_2603_vnum2 = 0;
_t___block_2608_cmp_yx = 0;
_t___block_2608_cmp_zx = 0;
_t___block_2608_cmp_zy = 0;
_t___block_2608_x_sel = 0;
_t___block_2608_y_sel = 0;
_t___block_2608_z_sel = 0;
_t___stage___block_2624_tex = 0;
_t___stage___block_2624_vnum0 = 0;
_t___stage___block_2624_vnum1 = 0;
_t___stage___block_2624_vnum2 = 0;
_t___block_2629_cmp_yx = 0;
_t___block_2629_cmp_zx = 0;
_t___block_2629_cmp_zy = 0;
_t___block_2629_x_sel = 0;
_t___block_2629_y_sel = 0;
_t___block_2629_z_sel = 0;
_t___stage___block_2645_tex = 0;
_t___stage___block_2645_vnum0 = 0;
_t___stage___block_2645_vnum1 = 0;
_t___stage___block_2645_vnum2 = 0;
_t___block_2650_cmp_yx = 0;
_t___block_2650_cmp_zx = 0;
_t___block_2650_cmp_zy = 0;
_t___block_2650_x_sel = 0;
_t___block_2650_y_sel = 0;
_t___block_2650_z_sel = 0;
_t___stage___block_2666_tex = 0;
_t___stage___block_2666_vnum0 = 0;
_t___stage___block_2666_vnum1 = 0;
_t___stage___block_2666_vnum2 = 0;
_t___block_2671_cmp_yx = 0;
_t___block_2671_cmp_zx = 0;
_t___block_2671_cmp_zy = 0;
_t___block_2671_x_sel = 0;
_t___block_2671_y_sel = 0;
_t___block_2671_z_sel = 0;
_t___stage___block_2687_tex = 0;
_t___stage___block_2687_vnum0 = 0;
_t___stage___block_2687_vnum1 = 0;
_t___stage___block_2687_vnum2 = 0;
_t___block_2692_cmp_yx = 0;
_t___block_2692_cmp_zx = 0;
_t___block_2692_cmp_zy = 0;
_t___block_2692_x_sel = 0;
_t___block_2692_y_sel = 0;
_t___block_2692_z_sel = 0;
_t___stage___block_2708_tex = 0;
_t___stage___block_2708_vnum0 = 0;
_t___stage___block_2708_vnum1 = 0;
_t___stage___block_2708_vnum2 = 0;
_t___block_2713_cmp_yx = 0;
_t___block_2713_cmp_zx = 0;
_t___block_2713_cmp_zy = 0;
_t___block_2713_x_sel = 0;
_t___block_2713_y_sel = 0;
_t___block_2713_z_sel = 0;
_t___stage___block_2729_fog = 0;
_t___stage___block_2729_light = 0;
_t___stage___block_2729_shade = 0;
_t___block_2731_clr_r = 0;
_t___block_2731_clr_g = 0;
_t___block_2731_clr_b = 0;
// _always_pre
(* full_case *)
case (_q__idx_fsm0)
1: begin
// _top
// __block_1
_d__idx_fsm0 = 2;
end
2: begin
// __while__block_2
if (1) begin
// __block_3
// __block_5
// --> pipeline __pip_5160_1 starts here
_t__1stdisable_fsm___pip_5160_1_0 = 0;
// __block_2738
// __block_2739
_d__idx_fsm0 = 2;
end else begin
// __block_4
// __block_2740
_d__idx_fsm0 = 0;
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
end
0: begin 
end
default: begin 
_d__idx_fsm0 = {2{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// ==== pipelines ====
// pipeline
// -------- stage 0
(* full_case *)
case (_q__idx_fsm___pip_5160_1_0)
1: begin
if (~_t__1stdisable_fsm___pip_5160_1_0) begin 
// __stage___block_6
// var inits
// --
_t___stage___block_6_vxsz = 1<<12;

_t___stage___block_6_view_x = (($signed(in_pix_x)-$signed(24'd320)));

_t___stage___block_6_view_y = (($signed(in_pix_y)-$signed(24'd240)));

_d_cos_addr0 = _q_frame>>1;

_d_sin_addr0 = _q_frame>>1;

_d_cos_addr1 = (_q_frame+(_q_frame<<1))>>3;

_d_sin_addr1 = (_q_frame+(_q_frame<<3))>>4;

// end of pipeline stage
_d__full_fsm___pip_5160_1_0 = 1;
end // 7
_d__idx_fsm___pip_5160_1_0 = _t__stall_fsm___pip_5160_1_0 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_0 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
if (_q__idx_fsm___pip_5160_1_0 == 1  ) begin
_d___pip_5160_1_0___stage___block_6_vxsz = _t___stage___block_6_vxsz;
end else begin
_d___pip_5160_1_0___stage___block_6_vxsz = _q___pip_5160_1_0___stage___block_6_vxsz;
end
if (_q__idx_fsm___pip_5160_1_0 == 1  ) begin
_d___pip_5160_1_0___stage___block_6_view_y = _t___stage___block_6_view_y;
end else begin
_d___pip_5160_1_0___stage___block_6_view_y = _q___pip_5160_1_0___stage___block_6_view_y;
end
if (_q__idx_fsm___pip_5160_1_0 == 1  ) begin
_d___pip_5160_1_0___stage___block_6_clr = _c___stage___block_6_clr;
end else begin
_d___pip_5160_1_0___stage___block_6_clr = _q___pip_5160_1_0___stage___block_6_clr;
end
if (_q__idx_fsm___pip_5160_1_0 == 1  ) begin
_d___pip_5160_1_0___stage___block_6_inside = _c___stage___block_6_inside;
end else begin
_d___pip_5160_1_0___stage___block_6_inside = _q___pip_5160_1_0___stage___block_6_inside;
end
if (_q__idx_fsm___pip_5160_1_0 == 1  ) begin
_d___pip_5160_1_0___stage___block_6_view_x = _t___stage___block_6_view_x;
end else begin
_d___pip_5160_1_0___stage___block_6_view_x = _q___pip_5160_1_0___stage___block_6_view_x;
end
if (_q__idx_fsm___pip_5160_1_0 == 1  ) begin
_d___pip_5160_1_0___stage___block_6_dist = _c___stage___block_6_dist;
end else begin
_d___pip_5160_1_0___stage___block_6_dist = _q___pip_5160_1_0___stage___block_6_dist;
end
if (_q__idx_fsm___pip_5160_1_0 == 1  ) begin
_d___pip_5160_1_0___stage___block_6_view_z = _c___stage___block_6_view_z;
end else begin
_d___pip_5160_1_0___stage___block_6_view_z = _q___pip_5160_1_0___stage___block_6_view_z;
end
// -------- stage 1
(* full_case *)
case (_q__idx_fsm___pip_5160_1_1)
1: begin
// __stage___block_7
_t___stage___block_7_cs0 = _w_mem_cos_rdata0;

_t___stage___block_7_ss0 = _w_mem_sin_rdata0;

_t___stage___block_7_cs1 = _w_mem_cos_rdata1;

_t___stage___block_7_ss1 = _w_mem_sin_rdata1;

// __block_8_imul_24_24
_t___stage___block_7_rot_x = _q___pip_5160_1_1___stage___block_6_view_x*_t___stage___block_7_cs1;

// __block_9
// __block_10_imul_24_24
_t___stage___block_7_rot_y = _q___pip_5160_1_1___stage___block_6_view_x*_t___stage___block_7_ss1;

// __block_11
// __block_12_imul_24_24
_t___block_11_yss = _q___pip_5160_1_1___stage___block_6_view_y*_t___stage___block_7_ss1;

// __block_13
// __block_14_imul_24_24
_t___block_11_ycs = _q___pip_5160_1_1___stage___block_6_view_y*_t___stage___block_7_cs1;

// __block_15
_d___pip_5160_1_1___stage___block_6_view_x = _t___stage___block_7_rot_x-_t___block_11_yss;

_d___pip_5160_1_1___stage___block_6_view_y = _t___stage___block_7_rot_y+_t___block_11_ycs;

// end of pipeline stage
_d__full_fsm___pip_5160_1_1 = 1;
_d__idx_fsm___pip_5160_1_1 = _t__stall_fsm___pip_5160_1_1 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_1 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
if (_q__idx_fsm___pip_5160_1_1 == 1  ) begin
_d___pip_5160_1_1___stage___block_7_ss0 = _t___stage___block_7_ss0;
end else begin
_d___pip_5160_1_1___stage___block_7_ss0 = _q___pip_5160_1_1___stage___block_7_ss0;
end
if (_q__idx_fsm___pip_5160_1_1 == 1  ) begin
_d___pip_5160_1_1___stage___block_7_cs0 = _t___stage___block_7_cs0;
end else begin
_d___pip_5160_1_1___stage___block_7_cs0 = _q___pip_5160_1_1___stage___block_7_cs0;
end
// -------- stage 2
(* full_case *)
case (_q__idx_fsm___pip_5160_1_2)
1: begin
// __stage___block_16
_d___pip_5160_1_2___stage___block_6_view_x = _q___pip_5160_1_2___stage___block_6_view_x>>>10;

_d___pip_5160_1_2___stage___block_6_view_y = _q___pip_5160_1_2___stage___block_6_view_y>>>10;

// end of pipeline stage
_d__full_fsm___pip_5160_1_2 = 1;
_d__idx_fsm___pip_5160_1_2 = _t__stall_fsm___pip_5160_1_2 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_2 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 3
(* full_case *)
case (_q__idx_fsm___pip_5160_1_3)
1: begin
// __stage___block_17
// __block_18_imul_24_24
_t___stage___block_17_xcs = _q___pip_5160_1_3___stage___block_6_view_x*_q___pip_5160_1_3___stage___block_7_cs0;

// __block_19
// __block_20_imul_24_24
_t___block_19_xss = _q___pip_5160_1_3___stage___block_6_view_x*_q___pip_5160_1_3___stage___block_7_ss0;

// __block_21
// __block_22_imul_24_24
_t___block_21_zcs = _q___pip_5160_1_3___stage___block_6_view_z*_q___pip_5160_1_3___stage___block_7_cs0;

// __block_23
// __block_24_imul_24_24
_t___block_23_zss = _q___pip_5160_1_3___stage___block_6_view_z*_q___pip_5160_1_3___stage___block_7_ss0;

// __block_25
_t___block_25_r_x_delta = (_t___stage___block_17_xcs-_t___block_23_zss);

_t___block_25_r_z_delta = (_t___block_19_xss+_t___block_21_zcs);

// end of pipeline stage
_d__full_fsm___pip_5160_1_3 = 1;
_d__idx_fsm___pip_5160_1_3 = _t__stall_fsm___pip_5160_1_3 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_3 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
if (_q__idx_fsm___pip_5160_1_3 == 1  ) begin
_d___pip_5160_1_3___block_25_r_z_delta = _t___block_25_r_z_delta;
end else begin
_d___pip_5160_1_3___block_25_r_z_delta = _q___pip_5160_1_3___block_25_r_z_delta;
end
if (_q__idx_fsm___pip_5160_1_3 == 1  ) begin
_d___pip_5160_1_3___block_25_r_x_delta = _t___block_25_r_x_delta;
end else begin
_d___pip_5160_1_3___block_25_r_x_delta = _q___pip_5160_1_3___block_25_r_x_delta;
end
// -------- stage 4
(* full_case *)
case (_q__idx_fsm___pip_5160_1_4)
1: begin
// __stage___block_26
_t___stage___block_26_rd_x = _q___pip_5160_1_4___block_25_r_x_delta>>>10;

_t___stage___block_26_rd_y = _q___pip_5160_1_4___stage___block_6_view_y;

_t___stage___block_26_rd_z = _q___pip_5160_1_4___block_25_r_z_delta>>>10;

_t___stage___block_26_s_x = _t___stage___block_26_rd_x<0 ? -1:1;

_t___stage___block_26_s_y = _t___stage___block_26_rd_y<0 ? -1:1;

_t___stage___block_26_s_z = _t___stage___block_26_rd_z<0 ? -1:1;

_d_invA_addr0 = _t___stage___block_26_rd_x<0 ? -_t___stage___block_26_rd_x:_t___stage___block_26_rd_x;

_d_invA_addr1 = _t___stage___block_26_rd_y<0 ? -_t___stage___block_26_rd_y:_t___stage___block_26_rd_y;

_d_invB_addr = _t___stage___block_26_rd_z<0 ? -_t___stage___block_26_rd_z:_t___stage___block_26_rd_z;

_t___stage___block_26_p_x = (68<<11);

_t___stage___block_26_p_y = (12<<11);

_t___stage___block_26_p_z = (_q_frame<<9);

_t___stage___block_26_v_x = _t___stage___block_26_p_x>>12;

_t___stage___block_26_v_y = _t___stage___block_26_p_y>>12;

_t___stage___block_26_v_z = _t___stage___block_26_p_z>>12;

_t___stage___block_26_brd_x = (_t___stage___block_26_p_x-(_t___stage___block_26_v_x<<12));

_t___stage___block_26_brd_y = (_t___stage___block_26_p_y-(_t___stage___block_26_v_y<<12));

_t___stage___block_26_brd_z = (_t___stage___block_26_p_z-(_t___stage___block_26_v_z<<12));

// end of pipeline stage
_d__full_fsm___pip_5160_1_4 = 1;
_d__idx_fsm___pip_5160_1_4 = _t__stall_fsm___pip_5160_1_4 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_4 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
if (_q__idx_fsm___pip_5160_1_4 == 1  ) begin
_d___pip_5160_1_4___stage___block_26_brd_x = _t___stage___block_26_brd_x;
end else begin
_d___pip_5160_1_4___stage___block_26_brd_x = _q___pip_5160_1_4___stage___block_26_brd_x;
end
if (_q__idx_fsm___pip_5160_1_4 == 1  ) begin
_d___pip_5160_1_4___stage___block_26_s_z = _t___stage___block_26_s_z;
end else begin
_d___pip_5160_1_4___stage___block_26_s_z = _q___pip_5160_1_4___stage___block_26_s_z;
end
if (_q__idx_fsm___pip_5160_1_4 == 1  ) begin
_d___pip_5160_1_4___stage___block_26_brd_y = _t___stage___block_26_brd_y;
end else begin
_d___pip_5160_1_4___stage___block_26_brd_y = _q___pip_5160_1_4___stage___block_26_brd_y;
end
if (_q__idx_fsm___pip_5160_1_4 == 1  ) begin
_d___pip_5160_1_4___stage___block_26_brd_z = _t___stage___block_26_brd_z;
end else begin
_d___pip_5160_1_4___stage___block_26_brd_z = _q___pip_5160_1_4___stage___block_26_brd_z;
end
if (_q__idx_fsm___pip_5160_1_4 == 1  ) begin
_d___pip_5160_1_4___stage___block_26_s_y = _t___stage___block_26_s_y;
end else begin
_d___pip_5160_1_4___stage___block_26_s_y = _q___pip_5160_1_4___stage___block_26_s_y;
end
if (_q__idx_fsm___pip_5160_1_4 == 1  ) begin
_d___pip_5160_1_4___stage___block_26_rd_x = _t___stage___block_26_rd_x;
end else begin
_d___pip_5160_1_4___stage___block_26_rd_x = _q___pip_5160_1_4___stage___block_26_rd_x;
end
if (_q__idx_fsm___pip_5160_1_4 == 1  ) begin
_d___pip_5160_1_4___stage___block_26_rd_y = _t___stage___block_26_rd_y;
end else begin
_d___pip_5160_1_4___stage___block_26_rd_y = _q___pip_5160_1_4___stage___block_26_rd_y;
end
if (_q__idx_fsm___pip_5160_1_4 == 1  ) begin
_d___pip_5160_1_4___stage___block_26_rd_z = _t___stage___block_26_rd_z;
end else begin
_d___pip_5160_1_4___stage___block_26_rd_z = _q___pip_5160_1_4___stage___block_26_rd_z;
end
if (_q__idx_fsm___pip_5160_1_4 == 1  ) begin
_d___pip_5160_1_4___stage___block_26_s_x = _t___stage___block_26_s_x;
end else begin
_d___pip_5160_1_4___stage___block_26_s_x = _q___pip_5160_1_4___stage___block_26_s_x;
end
if (_q__idx_fsm___pip_5160_1_4 == 1  ) begin
_d___pip_5160_1_4___stage___block_26_v_x = _t___stage___block_26_v_x;
end else begin
_d___pip_5160_1_4___stage___block_26_v_x = _q___pip_5160_1_4___stage___block_26_v_x;
end
if (_q__idx_fsm___pip_5160_1_4 == 1  ) begin
_d___pip_5160_1_4___stage___block_26_v_y = _t___stage___block_26_v_y;
end else begin
_d___pip_5160_1_4___stage___block_26_v_y = _q___pip_5160_1_4___stage___block_26_v_y;
end
if (_q__idx_fsm___pip_5160_1_4 == 1  ) begin
_d___pip_5160_1_4___stage___block_26_v_z = _t___stage___block_26_v_z;
end else begin
_d___pip_5160_1_4___stage___block_26_v_z = _q___pip_5160_1_4___stage___block_26_v_z;
end
// -------- stage 5
(* full_case *)
case (_q__idx_fsm___pip_5160_1_5)
1: begin
// __stage___block_27
_d___pip_5160_1_5___stage___block_26_brd_x = _q___pip_5160_1_5___stage___block_26_rd_x<0 ? (_q___pip_5160_1_5___stage___block_26_brd_x):(_q___pip_5160_1_5___stage___block_6_vxsz-_q___pip_5160_1_5___stage___block_26_brd_x);

_d___pip_5160_1_5___stage___block_26_brd_y = _q___pip_5160_1_5___stage___block_26_rd_y<0 ? (_q___pip_5160_1_5___stage___block_26_brd_y):(_q___pip_5160_1_5___stage___block_6_vxsz-_q___pip_5160_1_5___stage___block_26_brd_y);

_d___pip_5160_1_5___stage___block_26_brd_z = _q___pip_5160_1_5___stage___block_26_rd_z<0 ? (_q___pip_5160_1_5___stage___block_26_brd_z):(_q___pip_5160_1_5___stage___block_6_vxsz-_q___pip_5160_1_5___stage___block_26_brd_z);

// end of pipeline stage
_d__full_fsm___pip_5160_1_5 = 1;
_d__idx_fsm___pip_5160_1_5 = _t__stall_fsm___pip_5160_1_5 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_5 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 6
(* full_case *)
case (_q__idx_fsm___pip_5160_1_6)
1: begin
// __stage___block_28
_t___stage___block_28_inv_x = _w_mem_invA_rdata0;

_t___stage___block_28_inv_y = _w_mem_invA_rdata1;

_t___stage___block_28_inv_z = _w_mem_invB_rdata;

// __block_29_mul_14_18
_t___stage___block_28_tm_x_ = _q___pip_5160_1_6___stage___block_26_brd_x*_t___stage___block_28_inv_x;

// __block_30
// __block_31_mul_14_18
_t___stage___block_28_tm_y_ = _q___pip_5160_1_6___stage___block_26_brd_y*_t___stage___block_28_inv_y;

// __block_32
// __block_33_mul_14_18
_t___stage___block_28_tm_z_ = _q___pip_5160_1_6___stage___block_26_brd_z*_t___stage___block_28_inv_z;

// __block_34
_t___block_34_tm_x = _t___stage___block_28_tm_x_>>12;

_t___block_34_tm_y = _t___stage___block_28_tm_y_>>12;

_t___block_34_tm_z = _t___stage___block_28_tm_z_>>12;

// __block_35_mul_14_18
_t___block_34_dt_x_ = _q___pip_5160_1_6___stage___block_6_vxsz*_t___stage___block_28_inv_x;

// __block_36
// __block_37_mul_14_18
_t___block_34_dt_y_ = _q___pip_5160_1_6___stage___block_6_vxsz*_t___stage___block_28_inv_y;

// __block_38
// __block_39_mul_14_18
_t___block_34_dt_z_ = _q___pip_5160_1_6___stage___block_6_vxsz*_t___stage___block_28_inv_z;

// __block_40
_t___block_40_dt_x = (_t___block_34_dt_x_>>12)-1;

_t___block_40_dt_y = (_t___block_34_dt_y_>>12)-1;

_t___block_40_dt_z = (_t___block_34_dt_z_>>12)-1;

// end of pipeline stage
_d__full_fsm___pip_5160_1_6 = 1;
_d__idx_fsm___pip_5160_1_6 = _t__stall_fsm___pip_5160_1_6 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_6 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
if (_q__idx_fsm___pip_5160_1_6 == 1  ) begin
_d___pip_5160_1_6___block_40_dt_z = _t___block_40_dt_z;
end else begin
_d___pip_5160_1_6___block_40_dt_z = _q___pip_5160_1_6___block_40_dt_z;
end
if (_q__idx_fsm___pip_5160_1_6 == 1  ) begin
_d___pip_5160_1_6___block_40_dt_x = _t___block_40_dt_x;
end else begin
_d___pip_5160_1_6___block_40_dt_x = _q___pip_5160_1_6___block_40_dt_x;
end
if (_q__idx_fsm___pip_5160_1_6 == 1  ) begin
_d___pip_5160_1_6___block_34_tm_x = _t___block_34_tm_x;
end else begin
_d___pip_5160_1_6___block_34_tm_x = _q___pip_5160_1_6___block_34_tm_x;
end
if (_q__idx_fsm___pip_5160_1_6 == 1  ) begin
_d___pip_5160_1_6___block_34_tm_y = _t___block_34_tm_y;
end else begin
_d___pip_5160_1_6___block_34_tm_y = _q___pip_5160_1_6___block_34_tm_y;
end
if (_q__idx_fsm___pip_5160_1_6 == 1  ) begin
_d___pip_5160_1_6___block_40_dt_y = _t___block_40_dt_y;
end else begin
_d___pip_5160_1_6___block_40_dt_y = _q___pip_5160_1_6___block_40_dt_y;
end
if (_q__idx_fsm___pip_5160_1_6 == 1  ) begin
_d___pip_5160_1_6___block_34_tm_z = _t___block_34_tm_z;
end else begin
_d___pip_5160_1_6___block_34_tm_z = _q___pip_5160_1_6___block_34_tm_z;
end
// -------- stage 7
(* full_case *)
case (_q__idx_fsm___pip_5160_1_7)
1: begin
// __stage___block_41
_t___stage___block_41_tex = (_q___pip_5160_1_7___stage___block_26_v_x)^(_q___pip_5160_1_7___stage___block_26_v_y)^(_q___pip_5160_1_7___stage___block_26_v_z);

_t___stage___block_41_vnum0 = {_q___pip_5160_1_7___stage___block_26_v_z[0+:2],_q___pip_5160_1_7___stage___block_26_v_y[0+:2],_q___pip_5160_1_7___stage___block_26_v_x[0+:2]};

_t___stage___block_41_vnum1 = {_q___pip_5160_1_7___stage___block_26_v_z[2+:2],_q___pip_5160_1_7___stage___block_26_v_y[2+:2],_q___pip_5160_1_7___stage___block_26_v_x[2+:2]};

_t___stage___block_41_vnum2 = {_q___pip_5160_1_7___stage___block_26_v_z[4+:2],_q___pip_5160_1_7___stage___block_26_v_y[4+:2],_q___pip_5160_1_7___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_7___stage___block_6_inside&_w_tile[_t___stage___block_41_vnum0+:1]&_w_tile[_t___stage___block_41_vnum1+:1]&_w_tile[_t___stage___block_41_vnum2+:1]) begin
// __block_42
// __block_44
_d___pip_5160_1_7___stage___block_6_clr = _t___stage___block_41_tex;

_d___pip_5160_1_7___stage___block_6_dist = 0;

_d___pip_5160_1_7___stage___block_6_inside = 1;

// __block_45
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_43
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_46
_t___block_46_cmp_yx = _q___pip_5160_1_7___block_34_tm_y-_q___pip_5160_1_7___block_34_tm_x;

_t___block_46_cmp_zx = _q___pip_5160_1_7___block_34_tm_z-_q___pip_5160_1_7___block_34_tm_x;

_t___block_46_cmp_zy = _q___pip_5160_1_7___block_34_tm_z-_q___pip_5160_1_7___block_34_tm_y;

_t___block_46_x_sel = ~_t___block_46_cmp_yx[20+:1]&&~_t___block_46_cmp_zx[20+:1];

_t___block_46_y_sel = _t___block_46_cmp_yx[20+:1]&&~_t___block_46_cmp_zy[20+:1];

_t___block_46_z_sel = _t___block_46_cmp_zx[20+:1]&&_t___block_46_cmp_zy[20+:1];

if (_t___block_46_x_sel) begin
// __block_47
// __block_49
_d___pip_5160_1_7___stage___block_26_v_x = _q___pip_5160_1_7___stage___block_26_v_x+_q___pip_5160_1_7___stage___block_26_s_x;

_d___pip_5160_1_7___block_34_tm_x = _q___pip_5160_1_7___block_34_tm_x+_q___pip_5160_1_7___block_40_dt_x;

// __block_50
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_48
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_51
if (_t___block_46_y_sel) begin
// __block_52
// __block_54
_d___pip_5160_1_7___stage___block_26_v_y = _q___pip_5160_1_7___stage___block_26_v_y+_q___pip_5160_1_7___stage___block_26_s_y;

_d___pip_5160_1_7___block_34_tm_y = _q___pip_5160_1_7___block_34_tm_y+_q___pip_5160_1_7___block_40_dt_y;

// __block_55
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_53
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_56
if (_t___block_46_z_sel) begin
// __block_57
// __block_59
_d___pip_5160_1_7___stage___block_26_v_z = _q___pip_5160_1_7___stage___block_26_v_z+_q___pip_5160_1_7___stage___block_26_s_z;

_d___pip_5160_1_7___block_34_tm_z = _q___pip_5160_1_7___block_34_tm_z+_q___pip_5160_1_7___block_40_dt_z;

// __block_60
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_58
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_61
// end of pipeline stage
_d__full_fsm___pip_5160_1_7 = 1;
_d__idx_fsm___pip_5160_1_7 = _t__stall_fsm___pip_5160_1_7 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_7 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 8
(* full_case *)
case (_q__idx_fsm___pip_5160_1_8)
1: begin
// __stage___block_62
_t___stage___block_62_tex = (_q___pip_5160_1_8___stage___block_26_v_x)^(_q___pip_5160_1_8___stage___block_26_v_y)^(_q___pip_5160_1_8___stage___block_26_v_z);

_t___stage___block_62_vnum0 = {_q___pip_5160_1_8___stage___block_26_v_z[0+:2],_q___pip_5160_1_8___stage___block_26_v_y[0+:2],_q___pip_5160_1_8___stage___block_26_v_x[0+:2]};

_t___stage___block_62_vnum1 = {_q___pip_5160_1_8___stage___block_26_v_z[2+:2],_q___pip_5160_1_8___stage___block_26_v_y[2+:2],_q___pip_5160_1_8___stage___block_26_v_x[2+:2]};

_t___stage___block_62_vnum2 = {_q___pip_5160_1_8___stage___block_26_v_z[4+:2],_q___pip_5160_1_8___stage___block_26_v_y[4+:2],_q___pip_5160_1_8___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_8___stage___block_6_inside&_w_tile[_t___stage___block_62_vnum0+:1]&_w_tile[_t___stage___block_62_vnum1+:1]&_w_tile[_t___stage___block_62_vnum2+:1]) begin
// __block_63
// __block_65
_d___pip_5160_1_8___stage___block_6_clr = _t___stage___block_62_tex;

_d___pip_5160_1_8___stage___block_6_dist = 1;

_d___pip_5160_1_8___stage___block_6_inside = 1;

// __block_66
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_64
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_67
_t___block_67_cmp_yx = _q___pip_5160_1_8___block_34_tm_y-_q___pip_5160_1_8___block_34_tm_x;

_t___block_67_cmp_zx = _q___pip_5160_1_8___block_34_tm_z-_q___pip_5160_1_8___block_34_tm_x;

_t___block_67_cmp_zy = _q___pip_5160_1_8___block_34_tm_z-_q___pip_5160_1_8___block_34_tm_y;

_t___block_67_x_sel = ~_t___block_67_cmp_yx[20+:1]&&~_t___block_67_cmp_zx[20+:1];

_t___block_67_y_sel = _t___block_67_cmp_yx[20+:1]&&~_t___block_67_cmp_zy[20+:1];

_t___block_67_z_sel = _t___block_67_cmp_zx[20+:1]&&_t___block_67_cmp_zy[20+:1];

if (_t___block_67_x_sel) begin
// __block_68
// __block_70
_d___pip_5160_1_8___stage___block_26_v_x = _q___pip_5160_1_8___stage___block_26_v_x+_q___pip_5160_1_8___stage___block_26_s_x;

_d___pip_5160_1_8___block_34_tm_x = _q___pip_5160_1_8___block_34_tm_x+_q___pip_5160_1_8___block_40_dt_x;

// __block_71
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_69
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_72
if (_t___block_67_y_sel) begin
// __block_73
// __block_75
_d___pip_5160_1_8___stage___block_26_v_y = _q___pip_5160_1_8___stage___block_26_v_y+_q___pip_5160_1_8___stage___block_26_s_y;

_d___pip_5160_1_8___block_34_tm_y = _q___pip_5160_1_8___block_34_tm_y+_q___pip_5160_1_8___block_40_dt_y;

// __block_76
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_74
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_77
if (_t___block_67_z_sel) begin
// __block_78
// __block_80
_d___pip_5160_1_8___stage___block_26_v_z = _q___pip_5160_1_8___stage___block_26_v_z+_q___pip_5160_1_8___stage___block_26_s_z;

_d___pip_5160_1_8___block_34_tm_z = _q___pip_5160_1_8___block_34_tm_z+_q___pip_5160_1_8___block_40_dt_z;

// __block_81
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_79
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_82
// end of pipeline stage
_d__full_fsm___pip_5160_1_8 = 1;
_d__idx_fsm___pip_5160_1_8 = _t__stall_fsm___pip_5160_1_8 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_8 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 9
(* full_case *)
case (_q__idx_fsm___pip_5160_1_9)
1: begin
// __stage___block_83
_t___stage___block_83_tex = (_q___pip_5160_1_9___stage___block_26_v_x)^(_q___pip_5160_1_9___stage___block_26_v_y)^(_q___pip_5160_1_9___stage___block_26_v_z);

_t___stage___block_83_vnum0 = {_q___pip_5160_1_9___stage___block_26_v_z[0+:2],_q___pip_5160_1_9___stage___block_26_v_y[0+:2],_q___pip_5160_1_9___stage___block_26_v_x[0+:2]};

_t___stage___block_83_vnum1 = {_q___pip_5160_1_9___stage___block_26_v_z[2+:2],_q___pip_5160_1_9___stage___block_26_v_y[2+:2],_q___pip_5160_1_9___stage___block_26_v_x[2+:2]};

_t___stage___block_83_vnum2 = {_q___pip_5160_1_9___stage___block_26_v_z[4+:2],_q___pip_5160_1_9___stage___block_26_v_y[4+:2],_q___pip_5160_1_9___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_9___stage___block_6_inside&_w_tile[_t___stage___block_83_vnum0+:1]&_w_tile[_t___stage___block_83_vnum1+:1]&_w_tile[_t___stage___block_83_vnum2+:1]) begin
// __block_84
// __block_86
_d___pip_5160_1_9___stage___block_6_clr = _t___stage___block_83_tex;

_d___pip_5160_1_9___stage___block_6_dist = 3;

_d___pip_5160_1_9___stage___block_6_inside = 1;

// __block_87
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_85
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_88
_t___block_88_cmp_yx = _q___pip_5160_1_9___block_34_tm_y-_q___pip_5160_1_9___block_34_tm_x;

_t___block_88_cmp_zx = _q___pip_5160_1_9___block_34_tm_z-_q___pip_5160_1_9___block_34_tm_x;

_t___block_88_cmp_zy = _q___pip_5160_1_9___block_34_tm_z-_q___pip_5160_1_9___block_34_tm_y;

_t___block_88_x_sel = ~_t___block_88_cmp_yx[20+:1]&&~_t___block_88_cmp_zx[20+:1];

_t___block_88_y_sel = _t___block_88_cmp_yx[20+:1]&&~_t___block_88_cmp_zy[20+:1];

_t___block_88_z_sel = _t___block_88_cmp_zx[20+:1]&&_t___block_88_cmp_zy[20+:1];

if (_t___block_88_x_sel) begin
// __block_89
// __block_91
_d___pip_5160_1_9___stage___block_26_v_x = _q___pip_5160_1_9___stage___block_26_v_x+_q___pip_5160_1_9___stage___block_26_s_x;

_d___pip_5160_1_9___block_34_tm_x = _q___pip_5160_1_9___block_34_tm_x+_q___pip_5160_1_9___block_40_dt_x;

// __block_92
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_90
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_93
if (_t___block_88_y_sel) begin
// __block_94
// __block_96
_d___pip_5160_1_9___stage___block_26_v_y = _q___pip_5160_1_9___stage___block_26_v_y+_q___pip_5160_1_9___stage___block_26_s_y;

_d___pip_5160_1_9___block_34_tm_y = _q___pip_5160_1_9___block_34_tm_y+_q___pip_5160_1_9___block_40_dt_y;

// __block_97
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_95
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_98
if (_t___block_88_z_sel) begin
// __block_99
// __block_101
_d___pip_5160_1_9___stage___block_26_v_z = _q___pip_5160_1_9___stage___block_26_v_z+_q___pip_5160_1_9___stage___block_26_s_z;

_d___pip_5160_1_9___block_34_tm_z = _q___pip_5160_1_9___block_34_tm_z+_q___pip_5160_1_9___block_40_dt_z;

// __block_102
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_100
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_103
// end of pipeline stage
_d__full_fsm___pip_5160_1_9 = 1;
_d__idx_fsm___pip_5160_1_9 = _t__stall_fsm___pip_5160_1_9 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_9 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 10
(* full_case *)
case (_q__idx_fsm___pip_5160_1_10)
1: begin
// __stage___block_104
_t___stage___block_104_tex = (_q___pip_5160_1_10___stage___block_26_v_x)^(_q___pip_5160_1_10___stage___block_26_v_y)^(_q___pip_5160_1_10___stage___block_26_v_z);

_t___stage___block_104_vnum0 = {_q___pip_5160_1_10___stage___block_26_v_z[0+:2],_q___pip_5160_1_10___stage___block_26_v_y[0+:2],_q___pip_5160_1_10___stage___block_26_v_x[0+:2]};

_t___stage___block_104_vnum1 = {_q___pip_5160_1_10___stage___block_26_v_z[2+:2],_q___pip_5160_1_10___stage___block_26_v_y[2+:2],_q___pip_5160_1_10___stage___block_26_v_x[2+:2]};

_t___stage___block_104_vnum2 = {_q___pip_5160_1_10___stage___block_26_v_z[4+:2],_q___pip_5160_1_10___stage___block_26_v_y[4+:2],_q___pip_5160_1_10___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_10___stage___block_6_inside&_w_tile[_t___stage___block_104_vnum0+:1]&_w_tile[_t___stage___block_104_vnum1+:1]&_w_tile[_t___stage___block_104_vnum2+:1]) begin
// __block_105
// __block_107
_d___pip_5160_1_10___stage___block_6_clr = _t___stage___block_104_tex;

_d___pip_5160_1_10___stage___block_6_dist = 5;

_d___pip_5160_1_10___stage___block_6_inside = 1;

// __block_108
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_106
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_109
_t___block_109_cmp_yx = _q___pip_5160_1_10___block_34_tm_y-_q___pip_5160_1_10___block_34_tm_x;

_t___block_109_cmp_zx = _q___pip_5160_1_10___block_34_tm_z-_q___pip_5160_1_10___block_34_tm_x;

_t___block_109_cmp_zy = _q___pip_5160_1_10___block_34_tm_z-_q___pip_5160_1_10___block_34_tm_y;

_t___block_109_x_sel = ~_t___block_109_cmp_yx[20+:1]&&~_t___block_109_cmp_zx[20+:1];

_t___block_109_y_sel = _t___block_109_cmp_yx[20+:1]&&~_t___block_109_cmp_zy[20+:1];

_t___block_109_z_sel = _t___block_109_cmp_zx[20+:1]&&_t___block_109_cmp_zy[20+:1];

if (_t___block_109_x_sel) begin
// __block_110
// __block_112
_d___pip_5160_1_10___stage___block_26_v_x = _q___pip_5160_1_10___stage___block_26_v_x+_q___pip_5160_1_10___stage___block_26_s_x;

_d___pip_5160_1_10___block_34_tm_x = _q___pip_5160_1_10___block_34_tm_x+_q___pip_5160_1_10___block_40_dt_x;

// __block_113
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_111
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_114
if (_t___block_109_y_sel) begin
// __block_115
// __block_117
_d___pip_5160_1_10___stage___block_26_v_y = _q___pip_5160_1_10___stage___block_26_v_y+_q___pip_5160_1_10___stage___block_26_s_y;

_d___pip_5160_1_10___block_34_tm_y = _q___pip_5160_1_10___block_34_tm_y+_q___pip_5160_1_10___block_40_dt_y;

// __block_118
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_116
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_119
if (_t___block_109_z_sel) begin
// __block_120
// __block_122
_d___pip_5160_1_10___stage___block_26_v_z = _q___pip_5160_1_10___stage___block_26_v_z+_q___pip_5160_1_10___stage___block_26_s_z;

_d___pip_5160_1_10___block_34_tm_z = _q___pip_5160_1_10___block_34_tm_z+_q___pip_5160_1_10___block_40_dt_z;

// __block_123
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_121
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_124
// end of pipeline stage
_d__full_fsm___pip_5160_1_10 = 1;
_d__idx_fsm___pip_5160_1_10 = _t__stall_fsm___pip_5160_1_10 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_10 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 11
(* full_case *)
case (_q__idx_fsm___pip_5160_1_11)
1: begin
// __stage___block_125
_t___stage___block_125_tex = (_q___pip_5160_1_11___stage___block_26_v_x)^(_q___pip_5160_1_11___stage___block_26_v_y)^(_q___pip_5160_1_11___stage___block_26_v_z);

_t___stage___block_125_vnum0 = {_q___pip_5160_1_11___stage___block_26_v_z[0+:2],_q___pip_5160_1_11___stage___block_26_v_y[0+:2],_q___pip_5160_1_11___stage___block_26_v_x[0+:2]};

_t___stage___block_125_vnum1 = {_q___pip_5160_1_11___stage___block_26_v_z[2+:2],_q___pip_5160_1_11___stage___block_26_v_y[2+:2],_q___pip_5160_1_11___stage___block_26_v_x[2+:2]};

_t___stage___block_125_vnum2 = {_q___pip_5160_1_11___stage___block_26_v_z[4+:2],_q___pip_5160_1_11___stage___block_26_v_y[4+:2],_q___pip_5160_1_11___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_11___stage___block_6_inside&_w_tile[_t___stage___block_125_vnum0+:1]&_w_tile[_t___stage___block_125_vnum1+:1]&_w_tile[_t___stage___block_125_vnum2+:1]) begin
// __block_126
// __block_128
_d___pip_5160_1_11___stage___block_6_clr = _t___stage___block_125_tex;

_d___pip_5160_1_11___stage___block_6_dist = 7;

_d___pip_5160_1_11___stage___block_6_inside = 1;

// __block_129
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_127
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_130
_t___block_130_cmp_yx = _q___pip_5160_1_11___block_34_tm_y-_q___pip_5160_1_11___block_34_tm_x;

_t___block_130_cmp_zx = _q___pip_5160_1_11___block_34_tm_z-_q___pip_5160_1_11___block_34_tm_x;

_t___block_130_cmp_zy = _q___pip_5160_1_11___block_34_tm_z-_q___pip_5160_1_11___block_34_tm_y;

_t___block_130_x_sel = ~_t___block_130_cmp_yx[20+:1]&&~_t___block_130_cmp_zx[20+:1];

_t___block_130_y_sel = _t___block_130_cmp_yx[20+:1]&&~_t___block_130_cmp_zy[20+:1];

_t___block_130_z_sel = _t___block_130_cmp_zx[20+:1]&&_t___block_130_cmp_zy[20+:1];

if (_t___block_130_x_sel) begin
// __block_131
// __block_133
_d___pip_5160_1_11___stage___block_26_v_x = _q___pip_5160_1_11___stage___block_26_v_x+_q___pip_5160_1_11___stage___block_26_s_x;

_d___pip_5160_1_11___block_34_tm_x = _q___pip_5160_1_11___block_34_tm_x+_q___pip_5160_1_11___block_40_dt_x;

// __block_134
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_132
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_135
if (_t___block_130_y_sel) begin
// __block_136
// __block_138
_d___pip_5160_1_11___stage___block_26_v_y = _q___pip_5160_1_11___stage___block_26_v_y+_q___pip_5160_1_11___stage___block_26_s_y;

_d___pip_5160_1_11___block_34_tm_y = _q___pip_5160_1_11___block_34_tm_y+_q___pip_5160_1_11___block_40_dt_y;

// __block_139
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_137
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_140
if (_t___block_130_z_sel) begin
// __block_141
// __block_143
_d___pip_5160_1_11___stage___block_26_v_z = _q___pip_5160_1_11___stage___block_26_v_z+_q___pip_5160_1_11___stage___block_26_s_z;

_d___pip_5160_1_11___block_34_tm_z = _q___pip_5160_1_11___block_34_tm_z+_q___pip_5160_1_11___block_40_dt_z;

// __block_144
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_142
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_145
// end of pipeline stage
_d__full_fsm___pip_5160_1_11 = 1;
_d__idx_fsm___pip_5160_1_11 = _t__stall_fsm___pip_5160_1_11 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_11 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 12
(* full_case *)
case (_q__idx_fsm___pip_5160_1_12)
1: begin
// __stage___block_146
_t___stage___block_146_tex = (_q___pip_5160_1_12___stage___block_26_v_x)^(_q___pip_5160_1_12___stage___block_26_v_y)^(_q___pip_5160_1_12___stage___block_26_v_z);

_t___stage___block_146_vnum0 = {_q___pip_5160_1_12___stage___block_26_v_z[0+:2],_q___pip_5160_1_12___stage___block_26_v_y[0+:2],_q___pip_5160_1_12___stage___block_26_v_x[0+:2]};

_t___stage___block_146_vnum1 = {_q___pip_5160_1_12___stage___block_26_v_z[2+:2],_q___pip_5160_1_12___stage___block_26_v_y[2+:2],_q___pip_5160_1_12___stage___block_26_v_x[2+:2]};

_t___stage___block_146_vnum2 = {_q___pip_5160_1_12___stage___block_26_v_z[4+:2],_q___pip_5160_1_12___stage___block_26_v_y[4+:2],_q___pip_5160_1_12___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_12___stage___block_6_inside&_w_tile[_t___stage___block_146_vnum0+:1]&_w_tile[_t___stage___block_146_vnum1+:1]&_w_tile[_t___stage___block_146_vnum2+:1]) begin
// __block_147
// __block_149
_d___pip_5160_1_12___stage___block_6_clr = _t___stage___block_146_tex;

_d___pip_5160_1_12___stage___block_6_dist = 9;

_d___pip_5160_1_12___stage___block_6_inside = 1;

// __block_150
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_148
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_151
_t___block_151_cmp_yx = _q___pip_5160_1_12___block_34_tm_y-_q___pip_5160_1_12___block_34_tm_x;

_t___block_151_cmp_zx = _q___pip_5160_1_12___block_34_tm_z-_q___pip_5160_1_12___block_34_tm_x;

_t___block_151_cmp_zy = _q___pip_5160_1_12___block_34_tm_z-_q___pip_5160_1_12___block_34_tm_y;

_t___block_151_x_sel = ~_t___block_151_cmp_yx[20+:1]&&~_t___block_151_cmp_zx[20+:1];

_t___block_151_y_sel = _t___block_151_cmp_yx[20+:1]&&~_t___block_151_cmp_zy[20+:1];

_t___block_151_z_sel = _t___block_151_cmp_zx[20+:1]&&_t___block_151_cmp_zy[20+:1];

if (_t___block_151_x_sel) begin
// __block_152
// __block_154
_d___pip_5160_1_12___stage___block_26_v_x = _q___pip_5160_1_12___stage___block_26_v_x+_q___pip_5160_1_12___stage___block_26_s_x;

_d___pip_5160_1_12___block_34_tm_x = _q___pip_5160_1_12___block_34_tm_x+_q___pip_5160_1_12___block_40_dt_x;

// __block_155
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_153
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_156
if (_t___block_151_y_sel) begin
// __block_157
// __block_159
_d___pip_5160_1_12___stage___block_26_v_y = _q___pip_5160_1_12___stage___block_26_v_y+_q___pip_5160_1_12___stage___block_26_s_y;

_d___pip_5160_1_12___block_34_tm_y = _q___pip_5160_1_12___block_34_tm_y+_q___pip_5160_1_12___block_40_dt_y;

// __block_160
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_158
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_161
if (_t___block_151_z_sel) begin
// __block_162
// __block_164
_d___pip_5160_1_12___stage___block_26_v_z = _q___pip_5160_1_12___stage___block_26_v_z+_q___pip_5160_1_12___stage___block_26_s_z;

_d___pip_5160_1_12___block_34_tm_z = _q___pip_5160_1_12___block_34_tm_z+_q___pip_5160_1_12___block_40_dt_z;

// __block_165
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_163
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_166
// end of pipeline stage
_d__full_fsm___pip_5160_1_12 = 1;
_d__idx_fsm___pip_5160_1_12 = _t__stall_fsm___pip_5160_1_12 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_12 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 13
(* full_case *)
case (_q__idx_fsm___pip_5160_1_13)
1: begin
// __stage___block_167
_t___stage___block_167_tex = (_q___pip_5160_1_13___stage___block_26_v_x)^(_q___pip_5160_1_13___stage___block_26_v_y)^(_q___pip_5160_1_13___stage___block_26_v_z);

_t___stage___block_167_vnum0 = {_q___pip_5160_1_13___stage___block_26_v_z[0+:2],_q___pip_5160_1_13___stage___block_26_v_y[0+:2],_q___pip_5160_1_13___stage___block_26_v_x[0+:2]};

_t___stage___block_167_vnum1 = {_q___pip_5160_1_13___stage___block_26_v_z[2+:2],_q___pip_5160_1_13___stage___block_26_v_y[2+:2],_q___pip_5160_1_13___stage___block_26_v_x[2+:2]};

_t___stage___block_167_vnum2 = {_q___pip_5160_1_13___stage___block_26_v_z[4+:2],_q___pip_5160_1_13___stage___block_26_v_y[4+:2],_q___pip_5160_1_13___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_13___stage___block_6_inside&_w_tile[_t___stage___block_167_vnum0+:1]&_w_tile[_t___stage___block_167_vnum1+:1]&_w_tile[_t___stage___block_167_vnum2+:1]) begin
// __block_168
// __block_170
_d___pip_5160_1_13___stage___block_6_clr = _t___stage___block_167_tex;

_d___pip_5160_1_13___stage___block_6_dist = 11;

_d___pip_5160_1_13___stage___block_6_inside = 1;

// __block_171
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_169
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_172
_t___block_172_cmp_yx = _q___pip_5160_1_13___block_34_tm_y-_q___pip_5160_1_13___block_34_tm_x;

_t___block_172_cmp_zx = _q___pip_5160_1_13___block_34_tm_z-_q___pip_5160_1_13___block_34_tm_x;

_t___block_172_cmp_zy = _q___pip_5160_1_13___block_34_tm_z-_q___pip_5160_1_13___block_34_tm_y;

_t___block_172_x_sel = ~_t___block_172_cmp_yx[20+:1]&&~_t___block_172_cmp_zx[20+:1];

_t___block_172_y_sel = _t___block_172_cmp_yx[20+:1]&&~_t___block_172_cmp_zy[20+:1];

_t___block_172_z_sel = _t___block_172_cmp_zx[20+:1]&&_t___block_172_cmp_zy[20+:1];

if (_t___block_172_x_sel) begin
// __block_173
// __block_175
_d___pip_5160_1_13___stage___block_26_v_x = _q___pip_5160_1_13___stage___block_26_v_x+_q___pip_5160_1_13___stage___block_26_s_x;

_d___pip_5160_1_13___block_34_tm_x = _q___pip_5160_1_13___block_34_tm_x+_q___pip_5160_1_13___block_40_dt_x;

// __block_176
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_174
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_177
if (_t___block_172_y_sel) begin
// __block_178
// __block_180
_d___pip_5160_1_13___stage___block_26_v_y = _q___pip_5160_1_13___stage___block_26_v_y+_q___pip_5160_1_13___stage___block_26_s_y;

_d___pip_5160_1_13___block_34_tm_y = _q___pip_5160_1_13___block_34_tm_y+_q___pip_5160_1_13___block_40_dt_y;

// __block_181
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_179
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_182
if (_t___block_172_z_sel) begin
// __block_183
// __block_185
_d___pip_5160_1_13___stage___block_26_v_z = _q___pip_5160_1_13___stage___block_26_v_z+_q___pip_5160_1_13___stage___block_26_s_z;

_d___pip_5160_1_13___block_34_tm_z = _q___pip_5160_1_13___block_34_tm_z+_q___pip_5160_1_13___block_40_dt_z;

// __block_186
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_184
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_187
// end of pipeline stage
_d__full_fsm___pip_5160_1_13 = 1;
_d__idx_fsm___pip_5160_1_13 = _t__stall_fsm___pip_5160_1_13 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_13 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 14
(* full_case *)
case (_q__idx_fsm___pip_5160_1_14)
1: begin
// __stage___block_188
_t___stage___block_188_tex = (_q___pip_5160_1_14___stage___block_26_v_x)^(_q___pip_5160_1_14___stage___block_26_v_y)^(_q___pip_5160_1_14___stage___block_26_v_z);

_t___stage___block_188_vnum0 = {_q___pip_5160_1_14___stage___block_26_v_z[0+:2],_q___pip_5160_1_14___stage___block_26_v_y[0+:2],_q___pip_5160_1_14___stage___block_26_v_x[0+:2]};

_t___stage___block_188_vnum1 = {_q___pip_5160_1_14___stage___block_26_v_z[2+:2],_q___pip_5160_1_14___stage___block_26_v_y[2+:2],_q___pip_5160_1_14___stage___block_26_v_x[2+:2]};

_t___stage___block_188_vnum2 = {_q___pip_5160_1_14___stage___block_26_v_z[4+:2],_q___pip_5160_1_14___stage___block_26_v_y[4+:2],_q___pip_5160_1_14___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_14___stage___block_6_inside&_w_tile[_t___stage___block_188_vnum0+:1]&_w_tile[_t___stage___block_188_vnum1+:1]&_w_tile[_t___stage___block_188_vnum2+:1]) begin
// __block_189
// __block_191
_d___pip_5160_1_14___stage___block_6_clr = _t___stage___block_188_tex;

_d___pip_5160_1_14___stage___block_6_dist = 13;

_d___pip_5160_1_14___stage___block_6_inside = 1;

// __block_192
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_190
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_193
_t___block_193_cmp_yx = _q___pip_5160_1_14___block_34_tm_y-_q___pip_5160_1_14___block_34_tm_x;

_t___block_193_cmp_zx = _q___pip_5160_1_14___block_34_tm_z-_q___pip_5160_1_14___block_34_tm_x;

_t___block_193_cmp_zy = _q___pip_5160_1_14___block_34_tm_z-_q___pip_5160_1_14___block_34_tm_y;

_t___block_193_x_sel = ~_t___block_193_cmp_yx[20+:1]&&~_t___block_193_cmp_zx[20+:1];

_t___block_193_y_sel = _t___block_193_cmp_yx[20+:1]&&~_t___block_193_cmp_zy[20+:1];

_t___block_193_z_sel = _t___block_193_cmp_zx[20+:1]&&_t___block_193_cmp_zy[20+:1];

if (_t___block_193_x_sel) begin
// __block_194
// __block_196
_d___pip_5160_1_14___stage___block_26_v_x = _q___pip_5160_1_14___stage___block_26_v_x+_q___pip_5160_1_14___stage___block_26_s_x;

_d___pip_5160_1_14___block_34_tm_x = _q___pip_5160_1_14___block_34_tm_x+_q___pip_5160_1_14___block_40_dt_x;

// __block_197
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_195
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_198
if (_t___block_193_y_sel) begin
// __block_199
// __block_201
_d___pip_5160_1_14___stage___block_26_v_y = _q___pip_5160_1_14___stage___block_26_v_y+_q___pip_5160_1_14___stage___block_26_s_y;

_d___pip_5160_1_14___block_34_tm_y = _q___pip_5160_1_14___block_34_tm_y+_q___pip_5160_1_14___block_40_dt_y;

// __block_202
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_200
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_203
if (_t___block_193_z_sel) begin
// __block_204
// __block_206
_d___pip_5160_1_14___stage___block_26_v_z = _q___pip_5160_1_14___stage___block_26_v_z+_q___pip_5160_1_14___stage___block_26_s_z;

_d___pip_5160_1_14___block_34_tm_z = _q___pip_5160_1_14___block_34_tm_z+_q___pip_5160_1_14___block_40_dt_z;

// __block_207
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_205
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_208
// end of pipeline stage
_d__full_fsm___pip_5160_1_14 = 1;
_d__idx_fsm___pip_5160_1_14 = _t__stall_fsm___pip_5160_1_14 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_14 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 15
(* full_case *)
case (_q__idx_fsm___pip_5160_1_15)
1: begin
// __stage___block_209
_t___stage___block_209_tex = (_q___pip_5160_1_15___stage___block_26_v_x)^(_q___pip_5160_1_15___stage___block_26_v_y)^(_q___pip_5160_1_15___stage___block_26_v_z);

_t___stage___block_209_vnum0 = {_q___pip_5160_1_15___stage___block_26_v_z[0+:2],_q___pip_5160_1_15___stage___block_26_v_y[0+:2],_q___pip_5160_1_15___stage___block_26_v_x[0+:2]};

_t___stage___block_209_vnum1 = {_q___pip_5160_1_15___stage___block_26_v_z[2+:2],_q___pip_5160_1_15___stage___block_26_v_y[2+:2],_q___pip_5160_1_15___stage___block_26_v_x[2+:2]};

_t___stage___block_209_vnum2 = {_q___pip_5160_1_15___stage___block_26_v_z[4+:2],_q___pip_5160_1_15___stage___block_26_v_y[4+:2],_q___pip_5160_1_15___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_15___stage___block_6_inside&_w_tile[_t___stage___block_209_vnum0+:1]&_w_tile[_t___stage___block_209_vnum1+:1]&_w_tile[_t___stage___block_209_vnum2+:1]) begin
// __block_210
// __block_212
_d___pip_5160_1_15___stage___block_6_clr = _t___stage___block_209_tex;

_d___pip_5160_1_15___stage___block_6_dist = 14;

_d___pip_5160_1_15___stage___block_6_inside = 1;

// __block_213
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_211
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_214
_t___block_214_cmp_yx = _q___pip_5160_1_15___block_34_tm_y-_q___pip_5160_1_15___block_34_tm_x;

_t___block_214_cmp_zx = _q___pip_5160_1_15___block_34_tm_z-_q___pip_5160_1_15___block_34_tm_x;

_t___block_214_cmp_zy = _q___pip_5160_1_15___block_34_tm_z-_q___pip_5160_1_15___block_34_tm_y;

_t___block_214_x_sel = ~_t___block_214_cmp_yx[20+:1]&&~_t___block_214_cmp_zx[20+:1];

_t___block_214_y_sel = _t___block_214_cmp_yx[20+:1]&&~_t___block_214_cmp_zy[20+:1];

_t___block_214_z_sel = _t___block_214_cmp_zx[20+:1]&&_t___block_214_cmp_zy[20+:1];

if (_t___block_214_x_sel) begin
// __block_215
// __block_217
_d___pip_5160_1_15___stage___block_26_v_x = _q___pip_5160_1_15___stage___block_26_v_x+_q___pip_5160_1_15___stage___block_26_s_x;

_d___pip_5160_1_15___block_34_tm_x = _q___pip_5160_1_15___block_34_tm_x+_q___pip_5160_1_15___block_40_dt_x;

// __block_218
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_216
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_219
if (_t___block_214_y_sel) begin
// __block_220
// __block_222
_d___pip_5160_1_15___stage___block_26_v_y = _q___pip_5160_1_15___stage___block_26_v_y+_q___pip_5160_1_15___stage___block_26_s_y;

_d___pip_5160_1_15___block_34_tm_y = _q___pip_5160_1_15___block_34_tm_y+_q___pip_5160_1_15___block_40_dt_y;

// __block_223
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_221
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_224
if (_t___block_214_z_sel) begin
// __block_225
// __block_227
_d___pip_5160_1_15___stage___block_26_v_z = _q___pip_5160_1_15___stage___block_26_v_z+_q___pip_5160_1_15___stage___block_26_s_z;

_d___pip_5160_1_15___block_34_tm_z = _q___pip_5160_1_15___block_34_tm_z+_q___pip_5160_1_15___block_40_dt_z;

// __block_228
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_226
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_229
// end of pipeline stage
_d__full_fsm___pip_5160_1_15 = 1;
_d__idx_fsm___pip_5160_1_15 = _t__stall_fsm___pip_5160_1_15 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_15 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 16
(* full_case *)
case (_q__idx_fsm___pip_5160_1_16)
1: begin
// __stage___block_230
_t___stage___block_230_tex = (_q___pip_5160_1_16___stage___block_26_v_x)^(_q___pip_5160_1_16___stage___block_26_v_y)^(_q___pip_5160_1_16___stage___block_26_v_z);

_t___stage___block_230_vnum0 = {_q___pip_5160_1_16___stage___block_26_v_z[0+:2],_q___pip_5160_1_16___stage___block_26_v_y[0+:2],_q___pip_5160_1_16___stage___block_26_v_x[0+:2]};

_t___stage___block_230_vnum1 = {_q___pip_5160_1_16___stage___block_26_v_z[2+:2],_q___pip_5160_1_16___stage___block_26_v_y[2+:2],_q___pip_5160_1_16___stage___block_26_v_x[2+:2]};

_t___stage___block_230_vnum2 = {_q___pip_5160_1_16___stage___block_26_v_z[4+:2],_q___pip_5160_1_16___stage___block_26_v_y[4+:2],_q___pip_5160_1_16___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_16___stage___block_6_inside&_w_tile[_t___stage___block_230_vnum0+:1]&_w_tile[_t___stage___block_230_vnum1+:1]&_w_tile[_t___stage___block_230_vnum2+:1]) begin
// __block_231
// __block_233
_d___pip_5160_1_16___stage___block_6_clr = _t___stage___block_230_tex;

_d___pip_5160_1_16___stage___block_6_dist = 16;

_d___pip_5160_1_16___stage___block_6_inside = 1;

// __block_234
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_232
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_235
_t___block_235_cmp_yx = _q___pip_5160_1_16___block_34_tm_y-_q___pip_5160_1_16___block_34_tm_x;

_t___block_235_cmp_zx = _q___pip_5160_1_16___block_34_tm_z-_q___pip_5160_1_16___block_34_tm_x;

_t___block_235_cmp_zy = _q___pip_5160_1_16___block_34_tm_z-_q___pip_5160_1_16___block_34_tm_y;

_t___block_235_x_sel = ~_t___block_235_cmp_yx[20+:1]&&~_t___block_235_cmp_zx[20+:1];

_t___block_235_y_sel = _t___block_235_cmp_yx[20+:1]&&~_t___block_235_cmp_zy[20+:1];

_t___block_235_z_sel = _t___block_235_cmp_zx[20+:1]&&_t___block_235_cmp_zy[20+:1];

if (_t___block_235_x_sel) begin
// __block_236
// __block_238
_d___pip_5160_1_16___stage___block_26_v_x = _q___pip_5160_1_16___stage___block_26_v_x+_q___pip_5160_1_16___stage___block_26_s_x;

_d___pip_5160_1_16___block_34_tm_x = _q___pip_5160_1_16___block_34_tm_x+_q___pip_5160_1_16___block_40_dt_x;

// __block_239
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_237
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_240
if (_t___block_235_y_sel) begin
// __block_241
// __block_243
_d___pip_5160_1_16___stage___block_26_v_y = _q___pip_5160_1_16___stage___block_26_v_y+_q___pip_5160_1_16___stage___block_26_s_y;

_d___pip_5160_1_16___block_34_tm_y = _q___pip_5160_1_16___block_34_tm_y+_q___pip_5160_1_16___block_40_dt_y;

// __block_244
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_242
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_245
if (_t___block_235_z_sel) begin
// __block_246
// __block_248
_d___pip_5160_1_16___stage___block_26_v_z = _q___pip_5160_1_16___stage___block_26_v_z+_q___pip_5160_1_16___stage___block_26_s_z;

_d___pip_5160_1_16___block_34_tm_z = _q___pip_5160_1_16___block_34_tm_z+_q___pip_5160_1_16___block_40_dt_z;

// __block_249
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_247
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_250
// end of pipeline stage
_d__full_fsm___pip_5160_1_16 = 1;
_d__idx_fsm___pip_5160_1_16 = _t__stall_fsm___pip_5160_1_16 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_16 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 17
(* full_case *)
case (_q__idx_fsm___pip_5160_1_17)
1: begin
// __stage___block_251
_t___stage___block_251_tex = (_q___pip_5160_1_17___stage___block_26_v_x)^(_q___pip_5160_1_17___stage___block_26_v_y)^(_q___pip_5160_1_17___stage___block_26_v_z);

_t___stage___block_251_vnum0 = {_q___pip_5160_1_17___stage___block_26_v_z[0+:2],_q___pip_5160_1_17___stage___block_26_v_y[0+:2],_q___pip_5160_1_17___stage___block_26_v_x[0+:2]};

_t___stage___block_251_vnum1 = {_q___pip_5160_1_17___stage___block_26_v_z[2+:2],_q___pip_5160_1_17___stage___block_26_v_y[2+:2],_q___pip_5160_1_17___stage___block_26_v_x[2+:2]};

_t___stage___block_251_vnum2 = {_q___pip_5160_1_17___stage___block_26_v_z[4+:2],_q___pip_5160_1_17___stage___block_26_v_y[4+:2],_q___pip_5160_1_17___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_17___stage___block_6_inside&_w_tile[_t___stage___block_251_vnum0+:1]&_w_tile[_t___stage___block_251_vnum1+:1]&_w_tile[_t___stage___block_251_vnum2+:1]) begin
// __block_252
// __block_254
_d___pip_5160_1_17___stage___block_6_clr = _t___stage___block_251_tex;

_d___pip_5160_1_17___stage___block_6_dist = 18;

_d___pip_5160_1_17___stage___block_6_inside = 1;

// __block_255
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_253
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_256
_t___block_256_cmp_yx = _q___pip_5160_1_17___block_34_tm_y-_q___pip_5160_1_17___block_34_tm_x;

_t___block_256_cmp_zx = _q___pip_5160_1_17___block_34_tm_z-_q___pip_5160_1_17___block_34_tm_x;

_t___block_256_cmp_zy = _q___pip_5160_1_17___block_34_tm_z-_q___pip_5160_1_17___block_34_tm_y;

_t___block_256_x_sel = ~_t___block_256_cmp_yx[20+:1]&&~_t___block_256_cmp_zx[20+:1];

_t___block_256_y_sel = _t___block_256_cmp_yx[20+:1]&&~_t___block_256_cmp_zy[20+:1];

_t___block_256_z_sel = _t___block_256_cmp_zx[20+:1]&&_t___block_256_cmp_zy[20+:1];

if (_t___block_256_x_sel) begin
// __block_257
// __block_259
_d___pip_5160_1_17___stage___block_26_v_x = _q___pip_5160_1_17___stage___block_26_v_x+_q___pip_5160_1_17___stage___block_26_s_x;

_d___pip_5160_1_17___block_34_tm_x = _q___pip_5160_1_17___block_34_tm_x+_q___pip_5160_1_17___block_40_dt_x;

// __block_260
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_258
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_261
if (_t___block_256_y_sel) begin
// __block_262
// __block_264
_d___pip_5160_1_17___stage___block_26_v_y = _q___pip_5160_1_17___stage___block_26_v_y+_q___pip_5160_1_17___stage___block_26_s_y;

_d___pip_5160_1_17___block_34_tm_y = _q___pip_5160_1_17___block_34_tm_y+_q___pip_5160_1_17___block_40_dt_y;

// __block_265
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_263
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_266
if (_t___block_256_z_sel) begin
// __block_267
// __block_269
_d___pip_5160_1_17___stage___block_26_v_z = _q___pip_5160_1_17___stage___block_26_v_z+_q___pip_5160_1_17___stage___block_26_s_z;

_d___pip_5160_1_17___block_34_tm_z = _q___pip_5160_1_17___block_34_tm_z+_q___pip_5160_1_17___block_40_dt_z;

// __block_270
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_268
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_271
// end of pipeline stage
_d__full_fsm___pip_5160_1_17 = 1;
_d__idx_fsm___pip_5160_1_17 = _t__stall_fsm___pip_5160_1_17 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_17 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 18
(* full_case *)
case (_q__idx_fsm___pip_5160_1_18)
1: begin
// __stage___block_272
_t___stage___block_272_tex = (_q___pip_5160_1_18___stage___block_26_v_x)^(_q___pip_5160_1_18___stage___block_26_v_y)^(_q___pip_5160_1_18___stage___block_26_v_z);

_t___stage___block_272_vnum0 = {_q___pip_5160_1_18___stage___block_26_v_z[0+:2],_q___pip_5160_1_18___stage___block_26_v_y[0+:2],_q___pip_5160_1_18___stage___block_26_v_x[0+:2]};

_t___stage___block_272_vnum1 = {_q___pip_5160_1_18___stage___block_26_v_z[2+:2],_q___pip_5160_1_18___stage___block_26_v_y[2+:2],_q___pip_5160_1_18___stage___block_26_v_x[2+:2]};

_t___stage___block_272_vnum2 = {_q___pip_5160_1_18___stage___block_26_v_z[4+:2],_q___pip_5160_1_18___stage___block_26_v_y[4+:2],_q___pip_5160_1_18___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_18___stage___block_6_inside&_w_tile[_t___stage___block_272_vnum0+:1]&_w_tile[_t___stage___block_272_vnum1+:1]&_w_tile[_t___stage___block_272_vnum2+:1]) begin
// __block_273
// __block_275
_d___pip_5160_1_18___stage___block_6_clr = _t___stage___block_272_tex;

_d___pip_5160_1_18___stage___block_6_dist = 20;

_d___pip_5160_1_18___stage___block_6_inside = 1;

// __block_276
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_274
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_277
_t___block_277_cmp_yx = _q___pip_5160_1_18___block_34_tm_y-_q___pip_5160_1_18___block_34_tm_x;

_t___block_277_cmp_zx = _q___pip_5160_1_18___block_34_tm_z-_q___pip_5160_1_18___block_34_tm_x;

_t___block_277_cmp_zy = _q___pip_5160_1_18___block_34_tm_z-_q___pip_5160_1_18___block_34_tm_y;

_t___block_277_x_sel = ~_t___block_277_cmp_yx[20+:1]&&~_t___block_277_cmp_zx[20+:1];

_t___block_277_y_sel = _t___block_277_cmp_yx[20+:1]&&~_t___block_277_cmp_zy[20+:1];

_t___block_277_z_sel = _t___block_277_cmp_zx[20+:1]&&_t___block_277_cmp_zy[20+:1];

if (_t___block_277_x_sel) begin
// __block_278
// __block_280
_d___pip_5160_1_18___stage___block_26_v_x = _q___pip_5160_1_18___stage___block_26_v_x+_q___pip_5160_1_18___stage___block_26_s_x;

_d___pip_5160_1_18___block_34_tm_x = _q___pip_5160_1_18___block_34_tm_x+_q___pip_5160_1_18___block_40_dt_x;

// __block_281
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_279
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_282
if (_t___block_277_y_sel) begin
// __block_283
// __block_285
_d___pip_5160_1_18___stage___block_26_v_y = _q___pip_5160_1_18___stage___block_26_v_y+_q___pip_5160_1_18___stage___block_26_s_y;

_d___pip_5160_1_18___block_34_tm_y = _q___pip_5160_1_18___block_34_tm_y+_q___pip_5160_1_18___block_40_dt_y;

// __block_286
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_284
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_287
if (_t___block_277_z_sel) begin
// __block_288
// __block_290
_d___pip_5160_1_18___stage___block_26_v_z = _q___pip_5160_1_18___stage___block_26_v_z+_q___pip_5160_1_18___stage___block_26_s_z;

_d___pip_5160_1_18___block_34_tm_z = _q___pip_5160_1_18___block_34_tm_z+_q___pip_5160_1_18___block_40_dt_z;

// __block_291
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_289
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_292
// end of pipeline stage
_d__full_fsm___pip_5160_1_18 = 1;
_d__idx_fsm___pip_5160_1_18 = _t__stall_fsm___pip_5160_1_18 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_18 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 19
(* full_case *)
case (_q__idx_fsm___pip_5160_1_19)
1: begin
// __stage___block_293
_t___stage___block_293_tex = (_q___pip_5160_1_19___stage___block_26_v_x)^(_q___pip_5160_1_19___stage___block_26_v_y)^(_q___pip_5160_1_19___stage___block_26_v_z);

_t___stage___block_293_vnum0 = {_q___pip_5160_1_19___stage___block_26_v_z[0+:2],_q___pip_5160_1_19___stage___block_26_v_y[0+:2],_q___pip_5160_1_19___stage___block_26_v_x[0+:2]};

_t___stage___block_293_vnum1 = {_q___pip_5160_1_19___stage___block_26_v_z[2+:2],_q___pip_5160_1_19___stage___block_26_v_y[2+:2],_q___pip_5160_1_19___stage___block_26_v_x[2+:2]};

_t___stage___block_293_vnum2 = {_q___pip_5160_1_19___stage___block_26_v_z[4+:2],_q___pip_5160_1_19___stage___block_26_v_y[4+:2],_q___pip_5160_1_19___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_19___stage___block_6_inside&_w_tile[_t___stage___block_293_vnum0+:1]&_w_tile[_t___stage___block_293_vnum1+:1]&_w_tile[_t___stage___block_293_vnum2+:1]) begin
// __block_294
// __block_296
_d___pip_5160_1_19___stage___block_6_clr = _t___stage___block_293_tex;

_d___pip_5160_1_19___stage___block_6_dist = 22;

_d___pip_5160_1_19___stage___block_6_inside = 1;

// __block_297
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_295
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_298
_t___block_298_cmp_yx = _q___pip_5160_1_19___block_34_tm_y-_q___pip_5160_1_19___block_34_tm_x;

_t___block_298_cmp_zx = _q___pip_5160_1_19___block_34_tm_z-_q___pip_5160_1_19___block_34_tm_x;

_t___block_298_cmp_zy = _q___pip_5160_1_19___block_34_tm_z-_q___pip_5160_1_19___block_34_tm_y;

_t___block_298_x_sel = ~_t___block_298_cmp_yx[20+:1]&&~_t___block_298_cmp_zx[20+:1];

_t___block_298_y_sel = _t___block_298_cmp_yx[20+:1]&&~_t___block_298_cmp_zy[20+:1];

_t___block_298_z_sel = _t___block_298_cmp_zx[20+:1]&&_t___block_298_cmp_zy[20+:1];

if (_t___block_298_x_sel) begin
// __block_299
// __block_301
_d___pip_5160_1_19___stage___block_26_v_x = _q___pip_5160_1_19___stage___block_26_v_x+_q___pip_5160_1_19___stage___block_26_s_x;

_d___pip_5160_1_19___block_34_tm_x = _q___pip_5160_1_19___block_34_tm_x+_q___pip_5160_1_19___block_40_dt_x;

// __block_302
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_300
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_303
if (_t___block_298_y_sel) begin
// __block_304
// __block_306
_d___pip_5160_1_19___stage___block_26_v_y = _q___pip_5160_1_19___stage___block_26_v_y+_q___pip_5160_1_19___stage___block_26_s_y;

_d___pip_5160_1_19___block_34_tm_y = _q___pip_5160_1_19___block_34_tm_y+_q___pip_5160_1_19___block_40_dt_y;

// __block_307
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_305
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_308
if (_t___block_298_z_sel) begin
// __block_309
// __block_311
_d___pip_5160_1_19___stage___block_26_v_z = _q___pip_5160_1_19___stage___block_26_v_z+_q___pip_5160_1_19___stage___block_26_s_z;

_d___pip_5160_1_19___block_34_tm_z = _q___pip_5160_1_19___block_34_tm_z+_q___pip_5160_1_19___block_40_dt_z;

// __block_312
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_310
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_313
// end of pipeline stage
_d__full_fsm___pip_5160_1_19 = 1;
_d__idx_fsm___pip_5160_1_19 = _t__stall_fsm___pip_5160_1_19 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_19 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 20
(* full_case *)
case (_q__idx_fsm___pip_5160_1_20)
1: begin
// __stage___block_314
_t___stage___block_314_tex = (_q___pip_5160_1_20___stage___block_26_v_x)^(_q___pip_5160_1_20___stage___block_26_v_y)^(_q___pip_5160_1_20___stage___block_26_v_z);

_t___stage___block_314_vnum0 = {_q___pip_5160_1_20___stage___block_26_v_z[0+:2],_q___pip_5160_1_20___stage___block_26_v_y[0+:2],_q___pip_5160_1_20___stage___block_26_v_x[0+:2]};

_t___stage___block_314_vnum1 = {_q___pip_5160_1_20___stage___block_26_v_z[2+:2],_q___pip_5160_1_20___stage___block_26_v_y[2+:2],_q___pip_5160_1_20___stage___block_26_v_x[2+:2]};

_t___stage___block_314_vnum2 = {_q___pip_5160_1_20___stage___block_26_v_z[4+:2],_q___pip_5160_1_20___stage___block_26_v_y[4+:2],_q___pip_5160_1_20___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_20___stage___block_6_inside&_w_tile[_t___stage___block_314_vnum0+:1]&_w_tile[_t___stage___block_314_vnum1+:1]&_w_tile[_t___stage___block_314_vnum2+:1]) begin
// __block_315
// __block_317
_d___pip_5160_1_20___stage___block_6_clr = _t___stage___block_314_tex;

_d___pip_5160_1_20___stage___block_6_dist = 24;

_d___pip_5160_1_20___stage___block_6_inside = 1;

// __block_318
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_316
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_319
_t___block_319_cmp_yx = _q___pip_5160_1_20___block_34_tm_y-_q___pip_5160_1_20___block_34_tm_x;

_t___block_319_cmp_zx = _q___pip_5160_1_20___block_34_tm_z-_q___pip_5160_1_20___block_34_tm_x;

_t___block_319_cmp_zy = _q___pip_5160_1_20___block_34_tm_z-_q___pip_5160_1_20___block_34_tm_y;

_t___block_319_x_sel = ~_t___block_319_cmp_yx[20+:1]&&~_t___block_319_cmp_zx[20+:1];

_t___block_319_y_sel = _t___block_319_cmp_yx[20+:1]&&~_t___block_319_cmp_zy[20+:1];

_t___block_319_z_sel = _t___block_319_cmp_zx[20+:1]&&_t___block_319_cmp_zy[20+:1];

if (_t___block_319_x_sel) begin
// __block_320
// __block_322
_d___pip_5160_1_20___stage___block_26_v_x = _q___pip_5160_1_20___stage___block_26_v_x+_q___pip_5160_1_20___stage___block_26_s_x;

_d___pip_5160_1_20___block_34_tm_x = _q___pip_5160_1_20___block_34_tm_x+_q___pip_5160_1_20___block_40_dt_x;

// __block_323
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_321
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_324
if (_t___block_319_y_sel) begin
// __block_325
// __block_327
_d___pip_5160_1_20___stage___block_26_v_y = _q___pip_5160_1_20___stage___block_26_v_y+_q___pip_5160_1_20___stage___block_26_s_y;

_d___pip_5160_1_20___block_34_tm_y = _q___pip_5160_1_20___block_34_tm_y+_q___pip_5160_1_20___block_40_dt_y;

// __block_328
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_326
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_329
if (_t___block_319_z_sel) begin
// __block_330
// __block_332
_d___pip_5160_1_20___stage___block_26_v_z = _q___pip_5160_1_20___stage___block_26_v_z+_q___pip_5160_1_20___stage___block_26_s_z;

_d___pip_5160_1_20___block_34_tm_z = _q___pip_5160_1_20___block_34_tm_z+_q___pip_5160_1_20___block_40_dt_z;

// __block_333
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_331
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_334
// end of pipeline stage
_d__full_fsm___pip_5160_1_20 = 1;
_d__idx_fsm___pip_5160_1_20 = _t__stall_fsm___pip_5160_1_20 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_20 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 21
(* full_case *)
case (_q__idx_fsm___pip_5160_1_21)
1: begin
// __stage___block_335
_t___stage___block_335_tex = (_q___pip_5160_1_21___stage___block_26_v_x)^(_q___pip_5160_1_21___stage___block_26_v_y)^(_q___pip_5160_1_21___stage___block_26_v_z);

_t___stage___block_335_vnum0 = {_q___pip_5160_1_21___stage___block_26_v_z[0+:2],_q___pip_5160_1_21___stage___block_26_v_y[0+:2],_q___pip_5160_1_21___stage___block_26_v_x[0+:2]};

_t___stage___block_335_vnum1 = {_q___pip_5160_1_21___stage___block_26_v_z[2+:2],_q___pip_5160_1_21___stage___block_26_v_y[2+:2],_q___pip_5160_1_21___stage___block_26_v_x[2+:2]};

_t___stage___block_335_vnum2 = {_q___pip_5160_1_21___stage___block_26_v_z[4+:2],_q___pip_5160_1_21___stage___block_26_v_y[4+:2],_q___pip_5160_1_21___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_21___stage___block_6_inside&_w_tile[_t___stage___block_335_vnum0+:1]&_w_tile[_t___stage___block_335_vnum1+:1]&_w_tile[_t___stage___block_335_vnum2+:1]) begin
// __block_336
// __block_338
_d___pip_5160_1_21___stage___block_6_clr = _t___stage___block_335_tex;

_d___pip_5160_1_21___stage___block_6_dist = 26;

_d___pip_5160_1_21___stage___block_6_inside = 1;

// __block_339
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_337
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_340
_t___block_340_cmp_yx = _q___pip_5160_1_21___block_34_tm_y-_q___pip_5160_1_21___block_34_tm_x;

_t___block_340_cmp_zx = _q___pip_5160_1_21___block_34_tm_z-_q___pip_5160_1_21___block_34_tm_x;

_t___block_340_cmp_zy = _q___pip_5160_1_21___block_34_tm_z-_q___pip_5160_1_21___block_34_tm_y;

_t___block_340_x_sel = ~_t___block_340_cmp_yx[20+:1]&&~_t___block_340_cmp_zx[20+:1];

_t___block_340_y_sel = _t___block_340_cmp_yx[20+:1]&&~_t___block_340_cmp_zy[20+:1];

_t___block_340_z_sel = _t___block_340_cmp_zx[20+:1]&&_t___block_340_cmp_zy[20+:1];

if (_t___block_340_x_sel) begin
// __block_341
// __block_343
_d___pip_5160_1_21___stage___block_26_v_x = _q___pip_5160_1_21___stage___block_26_v_x+_q___pip_5160_1_21___stage___block_26_s_x;

_d___pip_5160_1_21___block_34_tm_x = _q___pip_5160_1_21___block_34_tm_x+_q___pip_5160_1_21___block_40_dt_x;

// __block_344
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_342
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_345
if (_t___block_340_y_sel) begin
// __block_346
// __block_348
_d___pip_5160_1_21___stage___block_26_v_y = _q___pip_5160_1_21___stage___block_26_v_y+_q___pip_5160_1_21___stage___block_26_s_y;

_d___pip_5160_1_21___block_34_tm_y = _q___pip_5160_1_21___block_34_tm_y+_q___pip_5160_1_21___block_40_dt_y;

// __block_349
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_347
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_350
if (_t___block_340_z_sel) begin
// __block_351
// __block_353
_d___pip_5160_1_21___stage___block_26_v_z = _q___pip_5160_1_21___stage___block_26_v_z+_q___pip_5160_1_21___stage___block_26_s_z;

_d___pip_5160_1_21___block_34_tm_z = _q___pip_5160_1_21___block_34_tm_z+_q___pip_5160_1_21___block_40_dt_z;

// __block_354
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_352
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_355
// end of pipeline stage
_d__full_fsm___pip_5160_1_21 = 1;
_d__idx_fsm___pip_5160_1_21 = _t__stall_fsm___pip_5160_1_21 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_21 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 22
(* full_case *)
case (_q__idx_fsm___pip_5160_1_22)
1: begin
// __stage___block_356
_t___stage___block_356_tex = (_q___pip_5160_1_22___stage___block_26_v_x)^(_q___pip_5160_1_22___stage___block_26_v_y)^(_q___pip_5160_1_22___stage___block_26_v_z);

_t___stage___block_356_vnum0 = {_q___pip_5160_1_22___stage___block_26_v_z[0+:2],_q___pip_5160_1_22___stage___block_26_v_y[0+:2],_q___pip_5160_1_22___stage___block_26_v_x[0+:2]};

_t___stage___block_356_vnum1 = {_q___pip_5160_1_22___stage___block_26_v_z[2+:2],_q___pip_5160_1_22___stage___block_26_v_y[2+:2],_q___pip_5160_1_22___stage___block_26_v_x[2+:2]};

_t___stage___block_356_vnum2 = {_q___pip_5160_1_22___stage___block_26_v_z[4+:2],_q___pip_5160_1_22___stage___block_26_v_y[4+:2],_q___pip_5160_1_22___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_22___stage___block_6_inside&_w_tile[_t___stage___block_356_vnum0+:1]&_w_tile[_t___stage___block_356_vnum1+:1]&_w_tile[_t___stage___block_356_vnum2+:1]) begin
// __block_357
// __block_359
_d___pip_5160_1_22___stage___block_6_clr = _t___stage___block_356_tex;

_d___pip_5160_1_22___stage___block_6_dist = 28;

_d___pip_5160_1_22___stage___block_6_inside = 1;

// __block_360
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_358
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_361
_t___block_361_cmp_yx = _q___pip_5160_1_22___block_34_tm_y-_q___pip_5160_1_22___block_34_tm_x;

_t___block_361_cmp_zx = _q___pip_5160_1_22___block_34_tm_z-_q___pip_5160_1_22___block_34_tm_x;

_t___block_361_cmp_zy = _q___pip_5160_1_22___block_34_tm_z-_q___pip_5160_1_22___block_34_tm_y;

_t___block_361_x_sel = ~_t___block_361_cmp_yx[20+:1]&&~_t___block_361_cmp_zx[20+:1];

_t___block_361_y_sel = _t___block_361_cmp_yx[20+:1]&&~_t___block_361_cmp_zy[20+:1];

_t___block_361_z_sel = _t___block_361_cmp_zx[20+:1]&&_t___block_361_cmp_zy[20+:1];

if (_t___block_361_x_sel) begin
// __block_362
// __block_364
_d___pip_5160_1_22___stage___block_26_v_x = _q___pip_5160_1_22___stage___block_26_v_x+_q___pip_5160_1_22___stage___block_26_s_x;

_d___pip_5160_1_22___block_34_tm_x = _q___pip_5160_1_22___block_34_tm_x+_q___pip_5160_1_22___block_40_dt_x;

// __block_365
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_363
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_366
if (_t___block_361_y_sel) begin
// __block_367
// __block_369
_d___pip_5160_1_22___stage___block_26_v_y = _q___pip_5160_1_22___stage___block_26_v_y+_q___pip_5160_1_22___stage___block_26_s_y;

_d___pip_5160_1_22___block_34_tm_y = _q___pip_5160_1_22___block_34_tm_y+_q___pip_5160_1_22___block_40_dt_y;

// __block_370
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_368
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_371
if (_t___block_361_z_sel) begin
// __block_372
// __block_374
_d___pip_5160_1_22___stage___block_26_v_z = _q___pip_5160_1_22___stage___block_26_v_z+_q___pip_5160_1_22___stage___block_26_s_z;

_d___pip_5160_1_22___block_34_tm_z = _q___pip_5160_1_22___block_34_tm_z+_q___pip_5160_1_22___block_40_dt_z;

// __block_375
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_373
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_376
// end of pipeline stage
_d__full_fsm___pip_5160_1_22 = 1;
_d__idx_fsm___pip_5160_1_22 = _t__stall_fsm___pip_5160_1_22 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_22 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 23
(* full_case *)
case (_q__idx_fsm___pip_5160_1_23)
1: begin
// __stage___block_377
_t___stage___block_377_tex = (_q___pip_5160_1_23___stage___block_26_v_x)^(_q___pip_5160_1_23___stage___block_26_v_y)^(_q___pip_5160_1_23___stage___block_26_v_z);

_t___stage___block_377_vnum0 = {_q___pip_5160_1_23___stage___block_26_v_z[0+:2],_q___pip_5160_1_23___stage___block_26_v_y[0+:2],_q___pip_5160_1_23___stage___block_26_v_x[0+:2]};

_t___stage___block_377_vnum1 = {_q___pip_5160_1_23___stage___block_26_v_z[2+:2],_q___pip_5160_1_23___stage___block_26_v_y[2+:2],_q___pip_5160_1_23___stage___block_26_v_x[2+:2]};

_t___stage___block_377_vnum2 = {_q___pip_5160_1_23___stage___block_26_v_z[4+:2],_q___pip_5160_1_23___stage___block_26_v_y[4+:2],_q___pip_5160_1_23___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_23___stage___block_6_inside&_w_tile[_t___stage___block_377_vnum0+:1]&_w_tile[_t___stage___block_377_vnum1+:1]&_w_tile[_t___stage___block_377_vnum2+:1]) begin
// __block_378
// __block_380
_d___pip_5160_1_23___stage___block_6_clr = _t___stage___block_377_tex;

_d___pip_5160_1_23___stage___block_6_dist = 29;

_d___pip_5160_1_23___stage___block_6_inside = 1;

// __block_381
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_379
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_382
_t___block_382_cmp_yx = _q___pip_5160_1_23___block_34_tm_y-_q___pip_5160_1_23___block_34_tm_x;

_t___block_382_cmp_zx = _q___pip_5160_1_23___block_34_tm_z-_q___pip_5160_1_23___block_34_tm_x;

_t___block_382_cmp_zy = _q___pip_5160_1_23___block_34_tm_z-_q___pip_5160_1_23___block_34_tm_y;

_t___block_382_x_sel = ~_t___block_382_cmp_yx[20+:1]&&~_t___block_382_cmp_zx[20+:1];

_t___block_382_y_sel = _t___block_382_cmp_yx[20+:1]&&~_t___block_382_cmp_zy[20+:1];

_t___block_382_z_sel = _t___block_382_cmp_zx[20+:1]&&_t___block_382_cmp_zy[20+:1];

if (_t___block_382_x_sel) begin
// __block_383
// __block_385
_d___pip_5160_1_23___stage___block_26_v_x = _q___pip_5160_1_23___stage___block_26_v_x+_q___pip_5160_1_23___stage___block_26_s_x;

_d___pip_5160_1_23___block_34_tm_x = _q___pip_5160_1_23___block_34_tm_x+_q___pip_5160_1_23___block_40_dt_x;

// __block_386
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_384
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_387
if (_t___block_382_y_sel) begin
// __block_388
// __block_390
_d___pip_5160_1_23___stage___block_26_v_y = _q___pip_5160_1_23___stage___block_26_v_y+_q___pip_5160_1_23___stage___block_26_s_y;

_d___pip_5160_1_23___block_34_tm_y = _q___pip_5160_1_23___block_34_tm_y+_q___pip_5160_1_23___block_40_dt_y;

// __block_391
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_389
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_392
if (_t___block_382_z_sel) begin
// __block_393
// __block_395
_d___pip_5160_1_23___stage___block_26_v_z = _q___pip_5160_1_23___stage___block_26_v_z+_q___pip_5160_1_23___stage___block_26_s_z;

_d___pip_5160_1_23___block_34_tm_z = _q___pip_5160_1_23___block_34_tm_z+_q___pip_5160_1_23___block_40_dt_z;

// __block_396
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_394
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_397
// end of pipeline stage
_d__full_fsm___pip_5160_1_23 = 1;
_d__idx_fsm___pip_5160_1_23 = _t__stall_fsm___pip_5160_1_23 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_23 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 24
(* full_case *)
case (_q__idx_fsm___pip_5160_1_24)
1: begin
// __stage___block_398
_t___stage___block_398_tex = (_q___pip_5160_1_24___stage___block_26_v_x)^(_q___pip_5160_1_24___stage___block_26_v_y)^(_q___pip_5160_1_24___stage___block_26_v_z);

_t___stage___block_398_vnum0 = {_q___pip_5160_1_24___stage___block_26_v_z[0+:2],_q___pip_5160_1_24___stage___block_26_v_y[0+:2],_q___pip_5160_1_24___stage___block_26_v_x[0+:2]};

_t___stage___block_398_vnum1 = {_q___pip_5160_1_24___stage___block_26_v_z[2+:2],_q___pip_5160_1_24___stage___block_26_v_y[2+:2],_q___pip_5160_1_24___stage___block_26_v_x[2+:2]};

_t___stage___block_398_vnum2 = {_q___pip_5160_1_24___stage___block_26_v_z[4+:2],_q___pip_5160_1_24___stage___block_26_v_y[4+:2],_q___pip_5160_1_24___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_24___stage___block_6_inside&_w_tile[_t___stage___block_398_vnum0+:1]&_w_tile[_t___stage___block_398_vnum1+:1]&_w_tile[_t___stage___block_398_vnum2+:1]) begin
// __block_399
// __block_401
_d___pip_5160_1_24___stage___block_6_clr = _t___stage___block_398_tex;

_d___pip_5160_1_24___stage___block_6_dist = 31;

_d___pip_5160_1_24___stage___block_6_inside = 1;

// __block_402
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_400
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_403
_t___block_403_cmp_yx = _q___pip_5160_1_24___block_34_tm_y-_q___pip_5160_1_24___block_34_tm_x;

_t___block_403_cmp_zx = _q___pip_5160_1_24___block_34_tm_z-_q___pip_5160_1_24___block_34_tm_x;

_t___block_403_cmp_zy = _q___pip_5160_1_24___block_34_tm_z-_q___pip_5160_1_24___block_34_tm_y;

_t___block_403_x_sel = ~_t___block_403_cmp_yx[20+:1]&&~_t___block_403_cmp_zx[20+:1];

_t___block_403_y_sel = _t___block_403_cmp_yx[20+:1]&&~_t___block_403_cmp_zy[20+:1];

_t___block_403_z_sel = _t___block_403_cmp_zx[20+:1]&&_t___block_403_cmp_zy[20+:1];

if (_t___block_403_x_sel) begin
// __block_404
// __block_406
_d___pip_5160_1_24___stage___block_26_v_x = _q___pip_5160_1_24___stage___block_26_v_x+_q___pip_5160_1_24___stage___block_26_s_x;

_d___pip_5160_1_24___block_34_tm_x = _q___pip_5160_1_24___block_34_tm_x+_q___pip_5160_1_24___block_40_dt_x;

// __block_407
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_405
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_408
if (_t___block_403_y_sel) begin
// __block_409
// __block_411
_d___pip_5160_1_24___stage___block_26_v_y = _q___pip_5160_1_24___stage___block_26_v_y+_q___pip_5160_1_24___stage___block_26_s_y;

_d___pip_5160_1_24___block_34_tm_y = _q___pip_5160_1_24___block_34_tm_y+_q___pip_5160_1_24___block_40_dt_y;

// __block_412
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_410
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_413
if (_t___block_403_z_sel) begin
// __block_414
// __block_416
_d___pip_5160_1_24___stage___block_26_v_z = _q___pip_5160_1_24___stage___block_26_v_z+_q___pip_5160_1_24___stage___block_26_s_z;

_d___pip_5160_1_24___block_34_tm_z = _q___pip_5160_1_24___block_34_tm_z+_q___pip_5160_1_24___block_40_dt_z;

// __block_417
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_415
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_418
// end of pipeline stage
_d__full_fsm___pip_5160_1_24 = 1;
_d__idx_fsm___pip_5160_1_24 = _t__stall_fsm___pip_5160_1_24 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_24 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 25
(* full_case *)
case (_q__idx_fsm___pip_5160_1_25)
1: begin
// __stage___block_419
_t___stage___block_419_tex = (_q___pip_5160_1_25___stage___block_26_v_x)^(_q___pip_5160_1_25___stage___block_26_v_y)^(_q___pip_5160_1_25___stage___block_26_v_z);

_t___stage___block_419_vnum0 = {_q___pip_5160_1_25___stage___block_26_v_z[0+:2],_q___pip_5160_1_25___stage___block_26_v_y[0+:2],_q___pip_5160_1_25___stage___block_26_v_x[0+:2]};

_t___stage___block_419_vnum1 = {_q___pip_5160_1_25___stage___block_26_v_z[2+:2],_q___pip_5160_1_25___stage___block_26_v_y[2+:2],_q___pip_5160_1_25___stage___block_26_v_x[2+:2]};

_t___stage___block_419_vnum2 = {_q___pip_5160_1_25___stage___block_26_v_z[4+:2],_q___pip_5160_1_25___stage___block_26_v_y[4+:2],_q___pip_5160_1_25___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_25___stage___block_6_inside&_w_tile[_t___stage___block_419_vnum0+:1]&_w_tile[_t___stage___block_419_vnum1+:1]&_w_tile[_t___stage___block_419_vnum2+:1]) begin
// __block_420
// __block_422
_d___pip_5160_1_25___stage___block_6_clr = _t___stage___block_419_tex;

_d___pip_5160_1_25___stage___block_6_dist = 33;

_d___pip_5160_1_25___stage___block_6_inside = 1;

// __block_423
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_421
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_424
_t___block_424_cmp_yx = _q___pip_5160_1_25___block_34_tm_y-_q___pip_5160_1_25___block_34_tm_x;

_t___block_424_cmp_zx = _q___pip_5160_1_25___block_34_tm_z-_q___pip_5160_1_25___block_34_tm_x;

_t___block_424_cmp_zy = _q___pip_5160_1_25___block_34_tm_z-_q___pip_5160_1_25___block_34_tm_y;

_t___block_424_x_sel = ~_t___block_424_cmp_yx[20+:1]&&~_t___block_424_cmp_zx[20+:1];

_t___block_424_y_sel = _t___block_424_cmp_yx[20+:1]&&~_t___block_424_cmp_zy[20+:1];

_t___block_424_z_sel = _t___block_424_cmp_zx[20+:1]&&_t___block_424_cmp_zy[20+:1];

if (_t___block_424_x_sel) begin
// __block_425
// __block_427
_d___pip_5160_1_25___stage___block_26_v_x = _q___pip_5160_1_25___stage___block_26_v_x+_q___pip_5160_1_25___stage___block_26_s_x;

_d___pip_5160_1_25___block_34_tm_x = _q___pip_5160_1_25___block_34_tm_x+_q___pip_5160_1_25___block_40_dt_x;

// __block_428
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_426
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_429
if (_t___block_424_y_sel) begin
// __block_430
// __block_432
_d___pip_5160_1_25___stage___block_26_v_y = _q___pip_5160_1_25___stage___block_26_v_y+_q___pip_5160_1_25___stage___block_26_s_y;

_d___pip_5160_1_25___block_34_tm_y = _q___pip_5160_1_25___block_34_tm_y+_q___pip_5160_1_25___block_40_dt_y;

// __block_433
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_431
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_434
if (_t___block_424_z_sel) begin
// __block_435
// __block_437
_d___pip_5160_1_25___stage___block_26_v_z = _q___pip_5160_1_25___stage___block_26_v_z+_q___pip_5160_1_25___stage___block_26_s_z;

_d___pip_5160_1_25___block_34_tm_z = _q___pip_5160_1_25___block_34_tm_z+_q___pip_5160_1_25___block_40_dt_z;

// __block_438
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_436
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_439
// end of pipeline stage
_d__full_fsm___pip_5160_1_25 = 1;
_d__idx_fsm___pip_5160_1_25 = _t__stall_fsm___pip_5160_1_25 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_25 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 26
(* full_case *)
case (_q__idx_fsm___pip_5160_1_26)
1: begin
// __stage___block_440
_t___stage___block_440_tex = (_q___pip_5160_1_26___stage___block_26_v_x)^(_q___pip_5160_1_26___stage___block_26_v_y)^(_q___pip_5160_1_26___stage___block_26_v_z);

_t___stage___block_440_vnum0 = {_q___pip_5160_1_26___stage___block_26_v_z[0+:2],_q___pip_5160_1_26___stage___block_26_v_y[0+:2],_q___pip_5160_1_26___stage___block_26_v_x[0+:2]};

_t___stage___block_440_vnum1 = {_q___pip_5160_1_26___stage___block_26_v_z[2+:2],_q___pip_5160_1_26___stage___block_26_v_y[2+:2],_q___pip_5160_1_26___stage___block_26_v_x[2+:2]};

_t___stage___block_440_vnum2 = {_q___pip_5160_1_26___stage___block_26_v_z[4+:2],_q___pip_5160_1_26___stage___block_26_v_y[4+:2],_q___pip_5160_1_26___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_26___stage___block_6_inside&_w_tile[_t___stage___block_440_vnum0+:1]&_w_tile[_t___stage___block_440_vnum1+:1]&_w_tile[_t___stage___block_440_vnum2+:1]) begin
// __block_441
// __block_443
_d___pip_5160_1_26___stage___block_6_clr = _t___stage___block_440_tex;

_d___pip_5160_1_26___stage___block_6_dist = 35;

_d___pip_5160_1_26___stage___block_6_inside = 1;

// __block_444
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_442
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_445
_t___block_445_cmp_yx = _q___pip_5160_1_26___block_34_tm_y-_q___pip_5160_1_26___block_34_tm_x;

_t___block_445_cmp_zx = _q___pip_5160_1_26___block_34_tm_z-_q___pip_5160_1_26___block_34_tm_x;

_t___block_445_cmp_zy = _q___pip_5160_1_26___block_34_tm_z-_q___pip_5160_1_26___block_34_tm_y;

_t___block_445_x_sel = ~_t___block_445_cmp_yx[20+:1]&&~_t___block_445_cmp_zx[20+:1];

_t___block_445_y_sel = _t___block_445_cmp_yx[20+:1]&&~_t___block_445_cmp_zy[20+:1];

_t___block_445_z_sel = _t___block_445_cmp_zx[20+:1]&&_t___block_445_cmp_zy[20+:1];

if (_t___block_445_x_sel) begin
// __block_446
// __block_448
_d___pip_5160_1_26___stage___block_26_v_x = _q___pip_5160_1_26___stage___block_26_v_x+_q___pip_5160_1_26___stage___block_26_s_x;

_d___pip_5160_1_26___block_34_tm_x = _q___pip_5160_1_26___block_34_tm_x+_q___pip_5160_1_26___block_40_dt_x;

// __block_449
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_447
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_450
if (_t___block_445_y_sel) begin
// __block_451
// __block_453
_d___pip_5160_1_26___stage___block_26_v_y = _q___pip_5160_1_26___stage___block_26_v_y+_q___pip_5160_1_26___stage___block_26_s_y;

_d___pip_5160_1_26___block_34_tm_y = _q___pip_5160_1_26___block_34_tm_y+_q___pip_5160_1_26___block_40_dt_y;

// __block_454
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_452
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_455
if (_t___block_445_z_sel) begin
// __block_456
// __block_458
_d___pip_5160_1_26___stage___block_26_v_z = _q___pip_5160_1_26___stage___block_26_v_z+_q___pip_5160_1_26___stage___block_26_s_z;

_d___pip_5160_1_26___block_34_tm_z = _q___pip_5160_1_26___block_34_tm_z+_q___pip_5160_1_26___block_40_dt_z;

// __block_459
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_457
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_460
// end of pipeline stage
_d__full_fsm___pip_5160_1_26 = 1;
_d__idx_fsm___pip_5160_1_26 = _t__stall_fsm___pip_5160_1_26 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_26 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 27
(* full_case *)
case (_q__idx_fsm___pip_5160_1_27)
1: begin
// __stage___block_461
_t___stage___block_461_tex = (_q___pip_5160_1_27___stage___block_26_v_x)^(_q___pip_5160_1_27___stage___block_26_v_y)^(_q___pip_5160_1_27___stage___block_26_v_z);

_t___stage___block_461_vnum0 = {_q___pip_5160_1_27___stage___block_26_v_z[0+:2],_q___pip_5160_1_27___stage___block_26_v_y[0+:2],_q___pip_5160_1_27___stage___block_26_v_x[0+:2]};

_t___stage___block_461_vnum1 = {_q___pip_5160_1_27___stage___block_26_v_z[2+:2],_q___pip_5160_1_27___stage___block_26_v_y[2+:2],_q___pip_5160_1_27___stage___block_26_v_x[2+:2]};

_t___stage___block_461_vnum2 = {_q___pip_5160_1_27___stage___block_26_v_z[4+:2],_q___pip_5160_1_27___stage___block_26_v_y[4+:2],_q___pip_5160_1_27___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_27___stage___block_6_inside&_w_tile[_t___stage___block_461_vnum0+:1]&_w_tile[_t___stage___block_461_vnum1+:1]&_w_tile[_t___stage___block_461_vnum2+:1]) begin
// __block_462
// __block_464
_d___pip_5160_1_27___stage___block_6_clr = _t___stage___block_461_tex;

_d___pip_5160_1_27___stage___block_6_dist = 37;

_d___pip_5160_1_27___stage___block_6_inside = 1;

// __block_465
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_463
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_466
_t___block_466_cmp_yx = _q___pip_5160_1_27___block_34_tm_y-_q___pip_5160_1_27___block_34_tm_x;

_t___block_466_cmp_zx = _q___pip_5160_1_27___block_34_tm_z-_q___pip_5160_1_27___block_34_tm_x;

_t___block_466_cmp_zy = _q___pip_5160_1_27___block_34_tm_z-_q___pip_5160_1_27___block_34_tm_y;

_t___block_466_x_sel = ~_t___block_466_cmp_yx[20+:1]&&~_t___block_466_cmp_zx[20+:1];

_t___block_466_y_sel = _t___block_466_cmp_yx[20+:1]&&~_t___block_466_cmp_zy[20+:1];

_t___block_466_z_sel = _t___block_466_cmp_zx[20+:1]&&_t___block_466_cmp_zy[20+:1];

if (_t___block_466_x_sel) begin
// __block_467
// __block_469
_d___pip_5160_1_27___stage___block_26_v_x = _q___pip_5160_1_27___stage___block_26_v_x+_q___pip_5160_1_27___stage___block_26_s_x;

_d___pip_5160_1_27___block_34_tm_x = _q___pip_5160_1_27___block_34_tm_x+_q___pip_5160_1_27___block_40_dt_x;

// __block_470
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_468
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_471
if (_t___block_466_y_sel) begin
// __block_472
// __block_474
_d___pip_5160_1_27___stage___block_26_v_y = _q___pip_5160_1_27___stage___block_26_v_y+_q___pip_5160_1_27___stage___block_26_s_y;

_d___pip_5160_1_27___block_34_tm_y = _q___pip_5160_1_27___block_34_tm_y+_q___pip_5160_1_27___block_40_dt_y;

// __block_475
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_473
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_476
if (_t___block_466_z_sel) begin
// __block_477
// __block_479
_d___pip_5160_1_27___stage___block_26_v_z = _q___pip_5160_1_27___stage___block_26_v_z+_q___pip_5160_1_27___stage___block_26_s_z;

_d___pip_5160_1_27___block_34_tm_z = _q___pip_5160_1_27___block_34_tm_z+_q___pip_5160_1_27___block_40_dt_z;

// __block_480
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_478
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_481
// end of pipeline stage
_d__full_fsm___pip_5160_1_27 = 1;
_d__idx_fsm___pip_5160_1_27 = _t__stall_fsm___pip_5160_1_27 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_27 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 28
(* full_case *)
case (_q__idx_fsm___pip_5160_1_28)
1: begin
// __stage___block_482
_t___stage___block_482_tex = (_q___pip_5160_1_28___stage___block_26_v_x)^(_q___pip_5160_1_28___stage___block_26_v_y)^(_q___pip_5160_1_28___stage___block_26_v_z);

_t___stage___block_482_vnum0 = {_q___pip_5160_1_28___stage___block_26_v_z[0+:2],_q___pip_5160_1_28___stage___block_26_v_y[0+:2],_q___pip_5160_1_28___stage___block_26_v_x[0+:2]};

_t___stage___block_482_vnum1 = {_q___pip_5160_1_28___stage___block_26_v_z[2+:2],_q___pip_5160_1_28___stage___block_26_v_y[2+:2],_q___pip_5160_1_28___stage___block_26_v_x[2+:2]};

_t___stage___block_482_vnum2 = {_q___pip_5160_1_28___stage___block_26_v_z[4+:2],_q___pip_5160_1_28___stage___block_26_v_y[4+:2],_q___pip_5160_1_28___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_28___stage___block_6_inside&_w_tile[_t___stage___block_482_vnum0+:1]&_w_tile[_t___stage___block_482_vnum1+:1]&_w_tile[_t___stage___block_482_vnum2+:1]) begin
// __block_483
// __block_485
_d___pip_5160_1_28___stage___block_6_clr = _t___stage___block_482_tex;

_d___pip_5160_1_28___stage___block_6_dist = 39;

_d___pip_5160_1_28___stage___block_6_inside = 1;

// __block_486
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_484
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_487
_t___block_487_cmp_yx = _q___pip_5160_1_28___block_34_tm_y-_q___pip_5160_1_28___block_34_tm_x;

_t___block_487_cmp_zx = _q___pip_5160_1_28___block_34_tm_z-_q___pip_5160_1_28___block_34_tm_x;

_t___block_487_cmp_zy = _q___pip_5160_1_28___block_34_tm_z-_q___pip_5160_1_28___block_34_tm_y;

_t___block_487_x_sel = ~_t___block_487_cmp_yx[20+:1]&&~_t___block_487_cmp_zx[20+:1];

_t___block_487_y_sel = _t___block_487_cmp_yx[20+:1]&&~_t___block_487_cmp_zy[20+:1];

_t___block_487_z_sel = _t___block_487_cmp_zx[20+:1]&&_t___block_487_cmp_zy[20+:1];

if (_t___block_487_x_sel) begin
// __block_488
// __block_490
_d___pip_5160_1_28___stage___block_26_v_x = _q___pip_5160_1_28___stage___block_26_v_x+_q___pip_5160_1_28___stage___block_26_s_x;

_d___pip_5160_1_28___block_34_tm_x = _q___pip_5160_1_28___block_34_tm_x+_q___pip_5160_1_28___block_40_dt_x;

// __block_491
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_489
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_492
if (_t___block_487_y_sel) begin
// __block_493
// __block_495
_d___pip_5160_1_28___stage___block_26_v_y = _q___pip_5160_1_28___stage___block_26_v_y+_q___pip_5160_1_28___stage___block_26_s_y;

_d___pip_5160_1_28___block_34_tm_y = _q___pip_5160_1_28___block_34_tm_y+_q___pip_5160_1_28___block_40_dt_y;

// __block_496
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_494
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_497
if (_t___block_487_z_sel) begin
// __block_498
// __block_500
_d___pip_5160_1_28___stage___block_26_v_z = _q___pip_5160_1_28___stage___block_26_v_z+_q___pip_5160_1_28___stage___block_26_s_z;

_d___pip_5160_1_28___block_34_tm_z = _q___pip_5160_1_28___block_34_tm_z+_q___pip_5160_1_28___block_40_dt_z;

// __block_501
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_499
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_502
// end of pipeline stage
_d__full_fsm___pip_5160_1_28 = 1;
_d__idx_fsm___pip_5160_1_28 = _t__stall_fsm___pip_5160_1_28 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_28 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 29
(* full_case *)
case (_q__idx_fsm___pip_5160_1_29)
1: begin
// __stage___block_503
_t___stage___block_503_tex = (_q___pip_5160_1_29___stage___block_26_v_x)^(_q___pip_5160_1_29___stage___block_26_v_y)^(_q___pip_5160_1_29___stage___block_26_v_z);

_t___stage___block_503_vnum0 = {_q___pip_5160_1_29___stage___block_26_v_z[0+:2],_q___pip_5160_1_29___stage___block_26_v_y[0+:2],_q___pip_5160_1_29___stage___block_26_v_x[0+:2]};

_t___stage___block_503_vnum1 = {_q___pip_5160_1_29___stage___block_26_v_z[2+:2],_q___pip_5160_1_29___stage___block_26_v_y[2+:2],_q___pip_5160_1_29___stage___block_26_v_x[2+:2]};

_t___stage___block_503_vnum2 = {_q___pip_5160_1_29___stage___block_26_v_z[4+:2],_q___pip_5160_1_29___stage___block_26_v_y[4+:2],_q___pip_5160_1_29___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_29___stage___block_6_inside&_w_tile[_t___stage___block_503_vnum0+:1]&_w_tile[_t___stage___block_503_vnum1+:1]&_w_tile[_t___stage___block_503_vnum2+:1]) begin
// __block_504
// __block_506
_d___pip_5160_1_29___stage___block_6_clr = _t___stage___block_503_tex;

_d___pip_5160_1_29___stage___block_6_dist = 41;

_d___pip_5160_1_29___stage___block_6_inside = 1;

// __block_507
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_505
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_508
_t___block_508_cmp_yx = _q___pip_5160_1_29___block_34_tm_y-_q___pip_5160_1_29___block_34_tm_x;

_t___block_508_cmp_zx = _q___pip_5160_1_29___block_34_tm_z-_q___pip_5160_1_29___block_34_tm_x;

_t___block_508_cmp_zy = _q___pip_5160_1_29___block_34_tm_z-_q___pip_5160_1_29___block_34_tm_y;

_t___block_508_x_sel = ~_t___block_508_cmp_yx[20+:1]&&~_t___block_508_cmp_zx[20+:1];

_t___block_508_y_sel = _t___block_508_cmp_yx[20+:1]&&~_t___block_508_cmp_zy[20+:1];

_t___block_508_z_sel = _t___block_508_cmp_zx[20+:1]&&_t___block_508_cmp_zy[20+:1];

if (_t___block_508_x_sel) begin
// __block_509
// __block_511
_d___pip_5160_1_29___stage___block_26_v_x = _q___pip_5160_1_29___stage___block_26_v_x+_q___pip_5160_1_29___stage___block_26_s_x;

_d___pip_5160_1_29___block_34_tm_x = _q___pip_5160_1_29___block_34_tm_x+_q___pip_5160_1_29___block_40_dt_x;

// __block_512
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_510
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_513
if (_t___block_508_y_sel) begin
// __block_514
// __block_516
_d___pip_5160_1_29___stage___block_26_v_y = _q___pip_5160_1_29___stage___block_26_v_y+_q___pip_5160_1_29___stage___block_26_s_y;

_d___pip_5160_1_29___block_34_tm_y = _q___pip_5160_1_29___block_34_tm_y+_q___pip_5160_1_29___block_40_dt_y;

// __block_517
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_515
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_518
if (_t___block_508_z_sel) begin
// __block_519
// __block_521
_d___pip_5160_1_29___stage___block_26_v_z = _q___pip_5160_1_29___stage___block_26_v_z+_q___pip_5160_1_29___stage___block_26_s_z;

_d___pip_5160_1_29___block_34_tm_z = _q___pip_5160_1_29___block_34_tm_z+_q___pip_5160_1_29___block_40_dt_z;

// __block_522
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_520
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_523
// end of pipeline stage
_d__full_fsm___pip_5160_1_29 = 1;
_d__idx_fsm___pip_5160_1_29 = _t__stall_fsm___pip_5160_1_29 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_29 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 30
(* full_case *)
case (_q__idx_fsm___pip_5160_1_30)
1: begin
// __stage___block_524
_t___stage___block_524_tex = (_q___pip_5160_1_30___stage___block_26_v_x)^(_q___pip_5160_1_30___stage___block_26_v_y)^(_q___pip_5160_1_30___stage___block_26_v_z);

_t___stage___block_524_vnum0 = {_q___pip_5160_1_30___stage___block_26_v_z[0+:2],_q___pip_5160_1_30___stage___block_26_v_y[0+:2],_q___pip_5160_1_30___stage___block_26_v_x[0+:2]};

_t___stage___block_524_vnum1 = {_q___pip_5160_1_30___stage___block_26_v_z[2+:2],_q___pip_5160_1_30___stage___block_26_v_y[2+:2],_q___pip_5160_1_30___stage___block_26_v_x[2+:2]};

_t___stage___block_524_vnum2 = {_q___pip_5160_1_30___stage___block_26_v_z[4+:2],_q___pip_5160_1_30___stage___block_26_v_y[4+:2],_q___pip_5160_1_30___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_30___stage___block_6_inside&_w_tile[_t___stage___block_524_vnum0+:1]&_w_tile[_t___stage___block_524_vnum1+:1]&_w_tile[_t___stage___block_524_vnum2+:1]) begin
// __block_525
// __block_527
_d___pip_5160_1_30___stage___block_6_clr = _t___stage___block_524_tex;

_d___pip_5160_1_30___stage___block_6_dist = 42;

_d___pip_5160_1_30___stage___block_6_inside = 1;

// __block_528
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_526
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_529
_t___block_529_cmp_yx = _q___pip_5160_1_30___block_34_tm_y-_q___pip_5160_1_30___block_34_tm_x;

_t___block_529_cmp_zx = _q___pip_5160_1_30___block_34_tm_z-_q___pip_5160_1_30___block_34_tm_x;

_t___block_529_cmp_zy = _q___pip_5160_1_30___block_34_tm_z-_q___pip_5160_1_30___block_34_tm_y;

_t___block_529_x_sel = ~_t___block_529_cmp_yx[20+:1]&&~_t___block_529_cmp_zx[20+:1];

_t___block_529_y_sel = _t___block_529_cmp_yx[20+:1]&&~_t___block_529_cmp_zy[20+:1];

_t___block_529_z_sel = _t___block_529_cmp_zx[20+:1]&&_t___block_529_cmp_zy[20+:1];

if (_t___block_529_x_sel) begin
// __block_530
// __block_532
_d___pip_5160_1_30___stage___block_26_v_x = _q___pip_5160_1_30___stage___block_26_v_x+_q___pip_5160_1_30___stage___block_26_s_x;

_d___pip_5160_1_30___block_34_tm_x = _q___pip_5160_1_30___block_34_tm_x+_q___pip_5160_1_30___block_40_dt_x;

// __block_533
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_531
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_534
if (_t___block_529_y_sel) begin
// __block_535
// __block_537
_d___pip_5160_1_30___stage___block_26_v_y = _q___pip_5160_1_30___stage___block_26_v_y+_q___pip_5160_1_30___stage___block_26_s_y;

_d___pip_5160_1_30___block_34_tm_y = _q___pip_5160_1_30___block_34_tm_y+_q___pip_5160_1_30___block_40_dt_y;

// __block_538
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_536
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_539
if (_t___block_529_z_sel) begin
// __block_540
// __block_542
_d___pip_5160_1_30___stage___block_26_v_z = _q___pip_5160_1_30___stage___block_26_v_z+_q___pip_5160_1_30___stage___block_26_s_z;

_d___pip_5160_1_30___block_34_tm_z = _q___pip_5160_1_30___block_34_tm_z+_q___pip_5160_1_30___block_40_dt_z;

// __block_543
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_541
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_544
// end of pipeline stage
_d__full_fsm___pip_5160_1_30 = 1;
_d__idx_fsm___pip_5160_1_30 = _t__stall_fsm___pip_5160_1_30 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_30 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 31
(* full_case *)
case (_q__idx_fsm___pip_5160_1_31)
1: begin
// __stage___block_545
_t___stage___block_545_tex = (_q___pip_5160_1_31___stage___block_26_v_x)^(_q___pip_5160_1_31___stage___block_26_v_y)^(_q___pip_5160_1_31___stage___block_26_v_z);

_t___stage___block_545_vnum0 = {_q___pip_5160_1_31___stage___block_26_v_z[0+:2],_q___pip_5160_1_31___stage___block_26_v_y[0+:2],_q___pip_5160_1_31___stage___block_26_v_x[0+:2]};

_t___stage___block_545_vnum1 = {_q___pip_5160_1_31___stage___block_26_v_z[2+:2],_q___pip_5160_1_31___stage___block_26_v_y[2+:2],_q___pip_5160_1_31___stage___block_26_v_x[2+:2]};

_t___stage___block_545_vnum2 = {_q___pip_5160_1_31___stage___block_26_v_z[4+:2],_q___pip_5160_1_31___stage___block_26_v_y[4+:2],_q___pip_5160_1_31___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_31___stage___block_6_inside&_w_tile[_t___stage___block_545_vnum0+:1]&_w_tile[_t___stage___block_545_vnum1+:1]&_w_tile[_t___stage___block_545_vnum2+:1]) begin
// __block_546
// __block_548
_d___pip_5160_1_31___stage___block_6_clr = _t___stage___block_545_tex;

_d___pip_5160_1_31___stage___block_6_dist = 44;

_d___pip_5160_1_31___stage___block_6_inside = 1;

// __block_549
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_547
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_550
_t___block_550_cmp_yx = _q___pip_5160_1_31___block_34_tm_y-_q___pip_5160_1_31___block_34_tm_x;

_t___block_550_cmp_zx = _q___pip_5160_1_31___block_34_tm_z-_q___pip_5160_1_31___block_34_tm_x;

_t___block_550_cmp_zy = _q___pip_5160_1_31___block_34_tm_z-_q___pip_5160_1_31___block_34_tm_y;

_t___block_550_x_sel = ~_t___block_550_cmp_yx[20+:1]&&~_t___block_550_cmp_zx[20+:1];

_t___block_550_y_sel = _t___block_550_cmp_yx[20+:1]&&~_t___block_550_cmp_zy[20+:1];

_t___block_550_z_sel = _t___block_550_cmp_zx[20+:1]&&_t___block_550_cmp_zy[20+:1];

if (_t___block_550_x_sel) begin
// __block_551
// __block_553
_d___pip_5160_1_31___stage___block_26_v_x = _q___pip_5160_1_31___stage___block_26_v_x+_q___pip_5160_1_31___stage___block_26_s_x;

_d___pip_5160_1_31___block_34_tm_x = _q___pip_5160_1_31___block_34_tm_x+_q___pip_5160_1_31___block_40_dt_x;

// __block_554
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_552
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_555
if (_t___block_550_y_sel) begin
// __block_556
// __block_558
_d___pip_5160_1_31___stage___block_26_v_y = _q___pip_5160_1_31___stage___block_26_v_y+_q___pip_5160_1_31___stage___block_26_s_y;

_d___pip_5160_1_31___block_34_tm_y = _q___pip_5160_1_31___block_34_tm_y+_q___pip_5160_1_31___block_40_dt_y;

// __block_559
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_557
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_560
if (_t___block_550_z_sel) begin
// __block_561
// __block_563
_d___pip_5160_1_31___stage___block_26_v_z = _q___pip_5160_1_31___stage___block_26_v_z+_q___pip_5160_1_31___stage___block_26_s_z;

_d___pip_5160_1_31___block_34_tm_z = _q___pip_5160_1_31___block_34_tm_z+_q___pip_5160_1_31___block_40_dt_z;

// __block_564
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_562
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_565
// end of pipeline stage
_d__full_fsm___pip_5160_1_31 = 1;
_d__idx_fsm___pip_5160_1_31 = _t__stall_fsm___pip_5160_1_31 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_31 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 32
(* full_case *)
case (_q__idx_fsm___pip_5160_1_32)
1: begin
// __stage___block_566
_t___stage___block_566_tex = (_q___pip_5160_1_32___stage___block_26_v_x)^(_q___pip_5160_1_32___stage___block_26_v_y)^(_q___pip_5160_1_32___stage___block_26_v_z);

_t___stage___block_566_vnum0 = {_q___pip_5160_1_32___stage___block_26_v_z[0+:2],_q___pip_5160_1_32___stage___block_26_v_y[0+:2],_q___pip_5160_1_32___stage___block_26_v_x[0+:2]};

_t___stage___block_566_vnum1 = {_q___pip_5160_1_32___stage___block_26_v_z[2+:2],_q___pip_5160_1_32___stage___block_26_v_y[2+:2],_q___pip_5160_1_32___stage___block_26_v_x[2+:2]};

_t___stage___block_566_vnum2 = {_q___pip_5160_1_32___stage___block_26_v_z[4+:2],_q___pip_5160_1_32___stage___block_26_v_y[4+:2],_q___pip_5160_1_32___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_32___stage___block_6_inside&_w_tile[_t___stage___block_566_vnum0+:1]&_w_tile[_t___stage___block_566_vnum1+:1]&_w_tile[_t___stage___block_566_vnum2+:1]) begin
// __block_567
// __block_569
_d___pip_5160_1_32___stage___block_6_clr = _t___stage___block_566_tex;

_d___pip_5160_1_32___stage___block_6_dist = 46;

_d___pip_5160_1_32___stage___block_6_inside = 1;

// __block_570
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_568
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_571
_t___block_571_cmp_yx = _q___pip_5160_1_32___block_34_tm_y-_q___pip_5160_1_32___block_34_tm_x;

_t___block_571_cmp_zx = _q___pip_5160_1_32___block_34_tm_z-_q___pip_5160_1_32___block_34_tm_x;

_t___block_571_cmp_zy = _q___pip_5160_1_32___block_34_tm_z-_q___pip_5160_1_32___block_34_tm_y;

_t___block_571_x_sel = ~_t___block_571_cmp_yx[20+:1]&&~_t___block_571_cmp_zx[20+:1];

_t___block_571_y_sel = _t___block_571_cmp_yx[20+:1]&&~_t___block_571_cmp_zy[20+:1];

_t___block_571_z_sel = _t___block_571_cmp_zx[20+:1]&&_t___block_571_cmp_zy[20+:1];

if (_t___block_571_x_sel) begin
// __block_572
// __block_574
_d___pip_5160_1_32___stage___block_26_v_x = _q___pip_5160_1_32___stage___block_26_v_x+_q___pip_5160_1_32___stage___block_26_s_x;

_d___pip_5160_1_32___block_34_tm_x = _q___pip_5160_1_32___block_34_tm_x+_q___pip_5160_1_32___block_40_dt_x;

// __block_575
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_573
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_576
if (_t___block_571_y_sel) begin
// __block_577
// __block_579
_d___pip_5160_1_32___stage___block_26_v_y = _q___pip_5160_1_32___stage___block_26_v_y+_q___pip_5160_1_32___stage___block_26_s_y;

_d___pip_5160_1_32___block_34_tm_y = _q___pip_5160_1_32___block_34_tm_y+_q___pip_5160_1_32___block_40_dt_y;

// __block_580
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_578
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_581
if (_t___block_571_z_sel) begin
// __block_582
// __block_584
_d___pip_5160_1_32___stage___block_26_v_z = _q___pip_5160_1_32___stage___block_26_v_z+_q___pip_5160_1_32___stage___block_26_s_z;

_d___pip_5160_1_32___block_34_tm_z = _q___pip_5160_1_32___block_34_tm_z+_q___pip_5160_1_32___block_40_dt_z;

// __block_585
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_583
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_586
// end of pipeline stage
_d__full_fsm___pip_5160_1_32 = 1;
_d__idx_fsm___pip_5160_1_32 = _t__stall_fsm___pip_5160_1_32 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_32 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 33
(* full_case *)
case (_q__idx_fsm___pip_5160_1_33)
1: begin
// __stage___block_587
_t___stage___block_587_tex = (_q___pip_5160_1_33___stage___block_26_v_x)^(_q___pip_5160_1_33___stage___block_26_v_y)^(_q___pip_5160_1_33___stage___block_26_v_z);

_t___stage___block_587_vnum0 = {_q___pip_5160_1_33___stage___block_26_v_z[0+:2],_q___pip_5160_1_33___stage___block_26_v_y[0+:2],_q___pip_5160_1_33___stage___block_26_v_x[0+:2]};

_t___stage___block_587_vnum1 = {_q___pip_5160_1_33___stage___block_26_v_z[2+:2],_q___pip_5160_1_33___stage___block_26_v_y[2+:2],_q___pip_5160_1_33___stage___block_26_v_x[2+:2]};

_t___stage___block_587_vnum2 = {_q___pip_5160_1_33___stage___block_26_v_z[4+:2],_q___pip_5160_1_33___stage___block_26_v_y[4+:2],_q___pip_5160_1_33___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_33___stage___block_6_inside&_w_tile[_t___stage___block_587_vnum0+:1]&_w_tile[_t___stage___block_587_vnum1+:1]&_w_tile[_t___stage___block_587_vnum2+:1]) begin
// __block_588
// __block_590
_d___pip_5160_1_33___stage___block_6_clr = _t___stage___block_587_tex;

_d___pip_5160_1_33___stage___block_6_dist = 48;

_d___pip_5160_1_33___stage___block_6_inside = 1;

// __block_591
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_589
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_592
_t___block_592_cmp_yx = _q___pip_5160_1_33___block_34_tm_y-_q___pip_5160_1_33___block_34_tm_x;

_t___block_592_cmp_zx = _q___pip_5160_1_33___block_34_tm_z-_q___pip_5160_1_33___block_34_tm_x;

_t___block_592_cmp_zy = _q___pip_5160_1_33___block_34_tm_z-_q___pip_5160_1_33___block_34_tm_y;

_t___block_592_x_sel = ~_t___block_592_cmp_yx[20+:1]&&~_t___block_592_cmp_zx[20+:1];

_t___block_592_y_sel = _t___block_592_cmp_yx[20+:1]&&~_t___block_592_cmp_zy[20+:1];

_t___block_592_z_sel = _t___block_592_cmp_zx[20+:1]&&_t___block_592_cmp_zy[20+:1];

if (_t___block_592_x_sel) begin
// __block_593
// __block_595
_d___pip_5160_1_33___stage___block_26_v_x = _q___pip_5160_1_33___stage___block_26_v_x+_q___pip_5160_1_33___stage___block_26_s_x;

_d___pip_5160_1_33___block_34_tm_x = _q___pip_5160_1_33___block_34_tm_x+_q___pip_5160_1_33___block_40_dt_x;

// __block_596
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_594
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_597
if (_t___block_592_y_sel) begin
// __block_598
// __block_600
_d___pip_5160_1_33___stage___block_26_v_y = _q___pip_5160_1_33___stage___block_26_v_y+_q___pip_5160_1_33___stage___block_26_s_y;

_d___pip_5160_1_33___block_34_tm_y = _q___pip_5160_1_33___block_34_tm_y+_q___pip_5160_1_33___block_40_dt_y;

// __block_601
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_599
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_602
if (_t___block_592_z_sel) begin
// __block_603
// __block_605
_d___pip_5160_1_33___stage___block_26_v_z = _q___pip_5160_1_33___stage___block_26_v_z+_q___pip_5160_1_33___stage___block_26_s_z;

_d___pip_5160_1_33___block_34_tm_z = _q___pip_5160_1_33___block_34_tm_z+_q___pip_5160_1_33___block_40_dt_z;

// __block_606
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_604
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_607
// end of pipeline stage
_d__full_fsm___pip_5160_1_33 = 1;
_d__idx_fsm___pip_5160_1_33 = _t__stall_fsm___pip_5160_1_33 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_33 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 34
(* full_case *)
case (_q__idx_fsm___pip_5160_1_34)
1: begin
// __stage___block_608
_t___stage___block_608_tex = (_q___pip_5160_1_34___stage___block_26_v_x)^(_q___pip_5160_1_34___stage___block_26_v_y)^(_q___pip_5160_1_34___stage___block_26_v_z);

_t___stage___block_608_vnum0 = {_q___pip_5160_1_34___stage___block_26_v_z[0+:2],_q___pip_5160_1_34___stage___block_26_v_y[0+:2],_q___pip_5160_1_34___stage___block_26_v_x[0+:2]};

_t___stage___block_608_vnum1 = {_q___pip_5160_1_34___stage___block_26_v_z[2+:2],_q___pip_5160_1_34___stage___block_26_v_y[2+:2],_q___pip_5160_1_34___stage___block_26_v_x[2+:2]};

_t___stage___block_608_vnum2 = {_q___pip_5160_1_34___stage___block_26_v_z[4+:2],_q___pip_5160_1_34___stage___block_26_v_y[4+:2],_q___pip_5160_1_34___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_34___stage___block_6_inside&_w_tile[_t___stage___block_608_vnum0+:1]&_w_tile[_t___stage___block_608_vnum1+:1]&_w_tile[_t___stage___block_608_vnum2+:1]) begin
// __block_609
// __block_611
_d___pip_5160_1_34___stage___block_6_clr = _t___stage___block_608_tex;

_d___pip_5160_1_34___stage___block_6_dist = 50;

_d___pip_5160_1_34___stage___block_6_inside = 1;

// __block_612
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_610
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_613
_t___block_613_cmp_yx = _q___pip_5160_1_34___block_34_tm_y-_q___pip_5160_1_34___block_34_tm_x;

_t___block_613_cmp_zx = _q___pip_5160_1_34___block_34_tm_z-_q___pip_5160_1_34___block_34_tm_x;

_t___block_613_cmp_zy = _q___pip_5160_1_34___block_34_tm_z-_q___pip_5160_1_34___block_34_tm_y;

_t___block_613_x_sel = ~_t___block_613_cmp_yx[20+:1]&&~_t___block_613_cmp_zx[20+:1];

_t___block_613_y_sel = _t___block_613_cmp_yx[20+:1]&&~_t___block_613_cmp_zy[20+:1];

_t___block_613_z_sel = _t___block_613_cmp_zx[20+:1]&&_t___block_613_cmp_zy[20+:1];

if (_t___block_613_x_sel) begin
// __block_614
// __block_616
_d___pip_5160_1_34___stage___block_26_v_x = _q___pip_5160_1_34___stage___block_26_v_x+_q___pip_5160_1_34___stage___block_26_s_x;

_d___pip_5160_1_34___block_34_tm_x = _q___pip_5160_1_34___block_34_tm_x+_q___pip_5160_1_34___block_40_dt_x;

// __block_617
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_615
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_618
if (_t___block_613_y_sel) begin
// __block_619
// __block_621
_d___pip_5160_1_34___stage___block_26_v_y = _q___pip_5160_1_34___stage___block_26_v_y+_q___pip_5160_1_34___stage___block_26_s_y;

_d___pip_5160_1_34___block_34_tm_y = _q___pip_5160_1_34___block_34_tm_y+_q___pip_5160_1_34___block_40_dt_y;

// __block_622
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_620
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_623
if (_t___block_613_z_sel) begin
// __block_624
// __block_626
_d___pip_5160_1_34___stage___block_26_v_z = _q___pip_5160_1_34___stage___block_26_v_z+_q___pip_5160_1_34___stage___block_26_s_z;

_d___pip_5160_1_34___block_34_tm_z = _q___pip_5160_1_34___block_34_tm_z+_q___pip_5160_1_34___block_40_dt_z;

// __block_627
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_625
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_628
// end of pipeline stage
_d__full_fsm___pip_5160_1_34 = 1;
_d__idx_fsm___pip_5160_1_34 = _t__stall_fsm___pip_5160_1_34 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_34 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 35
(* full_case *)
case (_q__idx_fsm___pip_5160_1_35)
1: begin
// __stage___block_629
_t___stage___block_629_tex = (_q___pip_5160_1_35___stage___block_26_v_x)^(_q___pip_5160_1_35___stage___block_26_v_y)^(_q___pip_5160_1_35___stage___block_26_v_z);

_t___stage___block_629_vnum0 = {_q___pip_5160_1_35___stage___block_26_v_z[0+:2],_q___pip_5160_1_35___stage___block_26_v_y[0+:2],_q___pip_5160_1_35___stage___block_26_v_x[0+:2]};

_t___stage___block_629_vnum1 = {_q___pip_5160_1_35___stage___block_26_v_z[2+:2],_q___pip_5160_1_35___stage___block_26_v_y[2+:2],_q___pip_5160_1_35___stage___block_26_v_x[2+:2]};

_t___stage___block_629_vnum2 = {_q___pip_5160_1_35___stage___block_26_v_z[4+:2],_q___pip_5160_1_35___stage___block_26_v_y[4+:2],_q___pip_5160_1_35___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_35___stage___block_6_inside&_w_tile[_t___stage___block_629_vnum0+:1]&_w_tile[_t___stage___block_629_vnum1+:1]&_w_tile[_t___stage___block_629_vnum2+:1]) begin
// __block_630
// __block_632
_d___pip_5160_1_35___stage___block_6_clr = _t___stage___block_629_tex;

_d___pip_5160_1_35___stage___block_6_dist = 52;

_d___pip_5160_1_35___stage___block_6_inside = 1;

// __block_633
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_631
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_634
_t___block_634_cmp_yx = _q___pip_5160_1_35___block_34_tm_y-_q___pip_5160_1_35___block_34_tm_x;

_t___block_634_cmp_zx = _q___pip_5160_1_35___block_34_tm_z-_q___pip_5160_1_35___block_34_tm_x;

_t___block_634_cmp_zy = _q___pip_5160_1_35___block_34_tm_z-_q___pip_5160_1_35___block_34_tm_y;

_t___block_634_x_sel = ~_t___block_634_cmp_yx[20+:1]&&~_t___block_634_cmp_zx[20+:1];

_t___block_634_y_sel = _t___block_634_cmp_yx[20+:1]&&~_t___block_634_cmp_zy[20+:1];

_t___block_634_z_sel = _t___block_634_cmp_zx[20+:1]&&_t___block_634_cmp_zy[20+:1];

if (_t___block_634_x_sel) begin
// __block_635
// __block_637
_d___pip_5160_1_35___stage___block_26_v_x = _q___pip_5160_1_35___stage___block_26_v_x+_q___pip_5160_1_35___stage___block_26_s_x;

_d___pip_5160_1_35___block_34_tm_x = _q___pip_5160_1_35___block_34_tm_x+_q___pip_5160_1_35___block_40_dt_x;

// __block_638
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_636
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_639
if (_t___block_634_y_sel) begin
// __block_640
// __block_642
_d___pip_5160_1_35___stage___block_26_v_y = _q___pip_5160_1_35___stage___block_26_v_y+_q___pip_5160_1_35___stage___block_26_s_y;

_d___pip_5160_1_35___block_34_tm_y = _q___pip_5160_1_35___block_34_tm_y+_q___pip_5160_1_35___block_40_dt_y;

// __block_643
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_641
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_644
if (_t___block_634_z_sel) begin
// __block_645
// __block_647
_d___pip_5160_1_35___stage___block_26_v_z = _q___pip_5160_1_35___stage___block_26_v_z+_q___pip_5160_1_35___stage___block_26_s_z;

_d___pip_5160_1_35___block_34_tm_z = _q___pip_5160_1_35___block_34_tm_z+_q___pip_5160_1_35___block_40_dt_z;

// __block_648
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_646
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_649
// end of pipeline stage
_d__full_fsm___pip_5160_1_35 = 1;
_d__idx_fsm___pip_5160_1_35 = _t__stall_fsm___pip_5160_1_35 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_35 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 36
(* full_case *)
case (_q__idx_fsm___pip_5160_1_36)
1: begin
// __stage___block_650
_t___stage___block_650_tex = (_q___pip_5160_1_36___stage___block_26_v_x)^(_q___pip_5160_1_36___stage___block_26_v_y)^(_q___pip_5160_1_36___stage___block_26_v_z);

_t___stage___block_650_vnum0 = {_q___pip_5160_1_36___stage___block_26_v_z[0+:2],_q___pip_5160_1_36___stage___block_26_v_y[0+:2],_q___pip_5160_1_36___stage___block_26_v_x[0+:2]};

_t___stage___block_650_vnum1 = {_q___pip_5160_1_36___stage___block_26_v_z[2+:2],_q___pip_5160_1_36___stage___block_26_v_y[2+:2],_q___pip_5160_1_36___stage___block_26_v_x[2+:2]};

_t___stage___block_650_vnum2 = {_q___pip_5160_1_36___stage___block_26_v_z[4+:2],_q___pip_5160_1_36___stage___block_26_v_y[4+:2],_q___pip_5160_1_36___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_36___stage___block_6_inside&_w_tile[_t___stage___block_650_vnum0+:1]&_w_tile[_t___stage___block_650_vnum1+:1]&_w_tile[_t___stage___block_650_vnum2+:1]) begin
// __block_651
// __block_653
_d___pip_5160_1_36___stage___block_6_clr = _t___stage___block_650_tex;

_d___pip_5160_1_36___stage___block_6_dist = 54;

_d___pip_5160_1_36___stage___block_6_inside = 1;

// __block_654
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_652
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_655
_t___block_655_cmp_yx = _q___pip_5160_1_36___block_34_tm_y-_q___pip_5160_1_36___block_34_tm_x;

_t___block_655_cmp_zx = _q___pip_5160_1_36___block_34_tm_z-_q___pip_5160_1_36___block_34_tm_x;

_t___block_655_cmp_zy = _q___pip_5160_1_36___block_34_tm_z-_q___pip_5160_1_36___block_34_tm_y;

_t___block_655_x_sel = ~_t___block_655_cmp_yx[20+:1]&&~_t___block_655_cmp_zx[20+:1];

_t___block_655_y_sel = _t___block_655_cmp_yx[20+:1]&&~_t___block_655_cmp_zy[20+:1];

_t___block_655_z_sel = _t___block_655_cmp_zx[20+:1]&&_t___block_655_cmp_zy[20+:1];

if (_t___block_655_x_sel) begin
// __block_656
// __block_658
_d___pip_5160_1_36___stage___block_26_v_x = _q___pip_5160_1_36___stage___block_26_v_x+_q___pip_5160_1_36___stage___block_26_s_x;

_d___pip_5160_1_36___block_34_tm_x = _q___pip_5160_1_36___block_34_tm_x+_q___pip_5160_1_36___block_40_dt_x;

// __block_659
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_657
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_660
if (_t___block_655_y_sel) begin
// __block_661
// __block_663
_d___pip_5160_1_36___stage___block_26_v_y = _q___pip_5160_1_36___stage___block_26_v_y+_q___pip_5160_1_36___stage___block_26_s_y;

_d___pip_5160_1_36___block_34_tm_y = _q___pip_5160_1_36___block_34_tm_y+_q___pip_5160_1_36___block_40_dt_y;

// __block_664
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_662
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_665
if (_t___block_655_z_sel) begin
// __block_666
// __block_668
_d___pip_5160_1_36___stage___block_26_v_z = _q___pip_5160_1_36___stage___block_26_v_z+_q___pip_5160_1_36___stage___block_26_s_z;

_d___pip_5160_1_36___block_34_tm_z = _q___pip_5160_1_36___block_34_tm_z+_q___pip_5160_1_36___block_40_dt_z;

// __block_669
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_667
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_670
// end of pipeline stage
_d__full_fsm___pip_5160_1_36 = 1;
_d__idx_fsm___pip_5160_1_36 = _t__stall_fsm___pip_5160_1_36 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_36 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 37
(* full_case *)
case (_q__idx_fsm___pip_5160_1_37)
1: begin
// __stage___block_671
_t___stage___block_671_tex = (_q___pip_5160_1_37___stage___block_26_v_x)^(_q___pip_5160_1_37___stage___block_26_v_y)^(_q___pip_5160_1_37___stage___block_26_v_z);

_t___stage___block_671_vnum0 = {_q___pip_5160_1_37___stage___block_26_v_z[0+:2],_q___pip_5160_1_37___stage___block_26_v_y[0+:2],_q___pip_5160_1_37___stage___block_26_v_x[0+:2]};

_t___stage___block_671_vnum1 = {_q___pip_5160_1_37___stage___block_26_v_z[2+:2],_q___pip_5160_1_37___stage___block_26_v_y[2+:2],_q___pip_5160_1_37___stage___block_26_v_x[2+:2]};

_t___stage___block_671_vnum2 = {_q___pip_5160_1_37___stage___block_26_v_z[4+:2],_q___pip_5160_1_37___stage___block_26_v_y[4+:2],_q___pip_5160_1_37___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_37___stage___block_6_inside&_w_tile[_t___stage___block_671_vnum0+:1]&_w_tile[_t___stage___block_671_vnum1+:1]&_w_tile[_t___stage___block_671_vnum2+:1]) begin
// __block_672
// __block_674
_d___pip_5160_1_37___stage___block_6_clr = _t___stage___block_671_tex;

_d___pip_5160_1_37___stage___block_6_dist = 56;

_d___pip_5160_1_37___stage___block_6_inside = 1;

// __block_675
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_673
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_676
_t___block_676_cmp_yx = _q___pip_5160_1_37___block_34_tm_y-_q___pip_5160_1_37___block_34_tm_x;

_t___block_676_cmp_zx = _q___pip_5160_1_37___block_34_tm_z-_q___pip_5160_1_37___block_34_tm_x;

_t___block_676_cmp_zy = _q___pip_5160_1_37___block_34_tm_z-_q___pip_5160_1_37___block_34_tm_y;

_t___block_676_x_sel = ~_t___block_676_cmp_yx[20+:1]&&~_t___block_676_cmp_zx[20+:1];

_t___block_676_y_sel = _t___block_676_cmp_yx[20+:1]&&~_t___block_676_cmp_zy[20+:1];

_t___block_676_z_sel = _t___block_676_cmp_zx[20+:1]&&_t___block_676_cmp_zy[20+:1];

if (_t___block_676_x_sel) begin
// __block_677
// __block_679
_d___pip_5160_1_37___stage___block_26_v_x = _q___pip_5160_1_37___stage___block_26_v_x+_q___pip_5160_1_37___stage___block_26_s_x;

_d___pip_5160_1_37___block_34_tm_x = _q___pip_5160_1_37___block_34_tm_x+_q___pip_5160_1_37___block_40_dt_x;

// __block_680
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_678
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_681
if (_t___block_676_y_sel) begin
// __block_682
// __block_684
_d___pip_5160_1_37___stage___block_26_v_y = _q___pip_5160_1_37___stage___block_26_v_y+_q___pip_5160_1_37___stage___block_26_s_y;

_d___pip_5160_1_37___block_34_tm_y = _q___pip_5160_1_37___block_34_tm_y+_q___pip_5160_1_37___block_40_dt_y;

// __block_685
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_683
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_686
if (_t___block_676_z_sel) begin
// __block_687
// __block_689
_d___pip_5160_1_37___stage___block_26_v_z = _q___pip_5160_1_37___stage___block_26_v_z+_q___pip_5160_1_37___stage___block_26_s_z;

_d___pip_5160_1_37___block_34_tm_z = _q___pip_5160_1_37___block_34_tm_z+_q___pip_5160_1_37___block_40_dt_z;

// __block_690
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_688
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_691
// end of pipeline stage
_d__full_fsm___pip_5160_1_37 = 1;
_d__idx_fsm___pip_5160_1_37 = _t__stall_fsm___pip_5160_1_37 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_37 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 38
(* full_case *)
case (_q__idx_fsm___pip_5160_1_38)
1: begin
// __stage___block_692
_t___stage___block_692_tex = (_q___pip_5160_1_38___stage___block_26_v_x)^(_q___pip_5160_1_38___stage___block_26_v_y)^(_q___pip_5160_1_38___stage___block_26_v_z);

_t___stage___block_692_vnum0 = {_q___pip_5160_1_38___stage___block_26_v_z[0+:2],_q___pip_5160_1_38___stage___block_26_v_y[0+:2],_q___pip_5160_1_38___stage___block_26_v_x[0+:2]};

_t___stage___block_692_vnum1 = {_q___pip_5160_1_38___stage___block_26_v_z[2+:2],_q___pip_5160_1_38___stage___block_26_v_y[2+:2],_q___pip_5160_1_38___stage___block_26_v_x[2+:2]};

_t___stage___block_692_vnum2 = {_q___pip_5160_1_38___stage___block_26_v_z[4+:2],_q___pip_5160_1_38___stage___block_26_v_y[4+:2],_q___pip_5160_1_38___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_38___stage___block_6_inside&_w_tile[_t___stage___block_692_vnum0+:1]&_w_tile[_t___stage___block_692_vnum1+:1]&_w_tile[_t___stage___block_692_vnum2+:1]) begin
// __block_693
// __block_695
_d___pip_5160_1_38___stage___block_6_clr = _t___stage___block_692_tex;

_d___pip_5160_1_38___stage___block_6_dist = 57;

_d___pip_5160_1_38___stage___block_6_inside = 1;

// __block_696
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_694
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_697
_t___block_697_cmp_yx = _q___pip_5160_1_38___block_34_tm_y-_q___pip_5160_1_38___block_34_tm_x;

_t___block_697_cmp_zx = _q___pip_5160_1_38___block_34_tm_z-_q___pip_5160_1_38___block_34_tm_x;

_t___block_697_cmp_zy = _q___pip_5160_1_38___block_34_tm_z-_q___pip_5160_1_38___block_34_tm_y;

_t___block_697_x_sel = ~_t___block_697_cmp_yx[20+:1]&&~_t___block_697_cmp_zx[20+:1];

_t___block_697_y_sel = _t___block_697_cmp_yx[20+:1]&&~_t___block_697_cmp_zy[20+:1];

_t___block_697_z_sel = _t___block_697_cmp_zx[20+:1]&&_t___block_697_cmp_zy[20+:1];

if (_t___block_697_x_sel) begin
// __block_698
// __block_700
_d___pip_5160_1_38___stage___block_26_v_x = _q___pip_5160_1_38___stage___block_26_v_x+_q___pip_5160_1_38___stage___block_26_s_x;

_d___pip_5160_1_38___block_34_tm_x = _q___pip_5160_1_38___block_34_tm_x+_q___pip_5160_1_38___block_40_dt_x;

// __block_701
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_699
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_702
if (_t___block_697_y_sel) begin
// __block_703
// __block_705
_d___pip_5160_1_38___stage___block_26_v_y = _q___pip_5160_1_38___stage___block_26_v_y+_q___pip_5160_1_38___stage___block_26_s_y;

_d___pip_5160_1_38___block_34_tm_y = _q___pip_5160_1_38___block_34_tm_y+_q___pip_5160_1_38___block_40_dt_y;

// __block_706
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_704
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_707
if (_t___block_697_z_sel) begin
// __block_708
// __block_710
_d___pip_5160_1_38___stage___block_26_v_z = _q___pip_5160_1_38___stage___block_26_v_z+_q___pip_5160_1_38___stage___block_26_s_z;

_d___pip_5160_1_38___block_34_tm_z = _q___pip_5160_1_38___block_34_tm_z+_q___pip_5160_1_38___block_40_dt_z;

// __block_711
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_709
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_712
// end of pipeline stage
_d__full_fsm___pip_5160_1_38 = 1;
_d__idx_fsm___pip_5160_1_38 = _t__stall_fsm___pip_5160_1_38 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_38 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 39
(* full_case *)
case (_q__idx_fsm___pip_5160_1_39)
1: begin
// __stage___block_713
_t___stage___block_713_tex = (_q___pip_5160_1_39___stage___block_26_v_x)^(_q___pip_5160_1_39___stage___block_26_v_y)^(_q___pip_5160_1_39___stage___block_26_v_z);

_t___stage___block_713_vnum0 = {_q___pip_5160_1_39___stage___block_26_v_z[0+:2],_q___pip_5160_1_39___stage___block_26_v_y[0+:2],_q___pip_5160_1_39___stage___block_26_v_x[0+:2]};

_t___stage___block_713_vnum1 = {_q___pip_5160_1_39___stage___block_26_v_z[2+:2],_q___pip_5160_1_39___stage___block_26_v_y[2+:2],_q___pip_5160_1_39___stage___block_26_v_x[2+:2]};

_t___stage___block_713_vnum2 = {_q___pip_5160_1_39___stage___block_26_v_z[4+:2],_q___pip_5160_1_39___stage___block_26_v_y[4+:2],_q___pip_5160_1_39___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_39___stage___block_6_inside&_w_tile[_t___stage___block_713_vnum0+:1]&_w_tile[_t___stage___block_713_vnum1+:1]&_w_tile[_t___stage___block_713_vnum2+:1]) begin
// __block_714
// __block_716
_d___pip_5160_1_39___stage___block_6_clr = _t___stage___block_713_tex;

_d___pip_5160_1_39___stage___block_6_dist = 59;

_d___pip_5160_1_39___stage___block_6_inside = 1;

// __block_717
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_715
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_718
_t___block_718_cmp_yx = _q___pip_5160_1_39___block_34_tm_y-_q___pip_5160_1_39___block_34_tm_x;

_t___block_718_cmp_zx = _q___pip_5160_1_39___block_34_tm_z-_q___pip_5160_1_39___block_34_tm_x;

_t___block_718_cmp_zy = _q___pip_5160_1_39___block_34_tm_z-_q___pip_5160_1_39___block_34_tm_y;

_t___block_718_x_sel = ~_t___block_718_cmp_yx[20+:1]&&~_t___block_718_cmp_zx[20+:1];

_t___block_718_y_sel = _t___block_718_cmp_yx[20+:1]&&~_t___block_718_cmp_zy[20+:1];

_t___block_718_z_sel = _t___block_718_cmp_zx[20+:1]&&_t___block_718_cmp_zy[20+:1];

if (_t___block_718_x_sel) begin
// __block_719
// __block_721
_d___pip_5160_1_39___stage___block_26_v_x = _q___pip_5160_1_39___stage___block_26_v_x+_q___pip_5160_1_39___stage___block_26_s_x;

_d___pip_5160_1_39___block_34_tm_x = _q___pip_5160_1_39___block_34_tm_x+_q___pip_5160_1_39___block_40_dt_x;

// __block_722
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_720
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_723
if (_t___block_718_y_sel) begin
// __block_724
// __block_726
_d___pip_5160_1_39___stage___block_26_v_y = _q___pip_5160_1_39___stage___block_26_v_y+_q___pip_5160_1_39___stage___block_26_s_y;

_d___pip_5160_1_39___block_34_tm_y = _q___pip_5160_1_39___block_34_tm_y+_q___pip_5160_1_39___block_40_dt_y;

// __block_727
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_725
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_728
if (_t___block_718_z_sel) begin
// __block_729
// __block_731
_d___pip_5160_1_39___stage___block_26_v_z = _q___pip_5160_1_39___stage___block_26_v_z+_q___pip_5160_1_39___stage___block_26_s_z;

_d___pip_5160_1_39___block_34_tm_z = _q___pip_5160_1_39___block_34_tm_z+_q___pip_5160_1_39___block_40_dt_z;

// __block_732
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_730
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_733
// end of pipeline stage
_d__full_fsm___pip_5160_1_39 = 1;
_d__idx_fsm___pip_5160_1_39 = _t__stall_fsm___pip_5160_1_39 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_39 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 40
(* full_case *)
case (_q__idx_fsm___pip_5160_1_40)
1: begin
// __stage___block_734
_t___stage___block_734_tex = (_q___pip_5160_1_40___stage___block_26_v_x)^(_q___pip_5160_1_40___stage___block_26_v_y)^(_q___pip_5160_1_40___stage___block_26_v_z);

_t___stage___block_734_vnum0 = {_q___pip_5160_1_40___stage___block_26_v_z[0+:2],_q___pip_5160_1_40___stage___block_26_v_y[0+:2],_q___pip_5160_1_40___stage___block_26_v_x[0+:2]};

_t___stage___block_734_vnum1 = {_q___pip_5160_1_40___stage___block_26_v_z[2+:2],_q___pip_5160_1_40___stage___block_26_v_y[2+:2],_q___pip_5160_1_40___stage___block_26_v_x[2+:2]};

_t___stage___block_734_vnum2 = {_q___pip_5160_1_40___stage___block_26_v_z[4+:2],_q___pip_5160_1_40___stage___block_26_v_y[4+:2],_q___pip_5160_1_40___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_40___stage___block_6_inside&_w_tile[_t___stage___block_734_vnum0+:1]&_w_tile[_t___stage___block_734_vnum1+:1]&_w_tile[_t___stage___block_734_vnum2+:1]) begin
// __block_735
// __block_737
_d___pip_5160_1_40___stage___block_6_clr = _t___stage___block_734_tex;

_d___pip_5160_1_40___stage___block_6_dist = 61;

_d___pip_5160_1_40___stage___block_6_inside = 1;

// __block_738
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_736
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_739
_t___block_739_cmp_yx = _q___pip_5160_1_40___block_34_tm_y-_q___pip_5160_1_40___block_34_tm_x;

_t___block_739_cmp_zx = _q___pip_5160_1_40___block_34_tm_z-_q___pip_5160_1_40___block_34_tm_x;

_t___block_739_cmp_zy = _q___pip_5160_1_40___block_34_tm_z-_q___pip_5160_1_40___block_34_tm_y;

_t___block_739_x_sel = ~_t___block_739_cmp_yx[20+:1]&&~_t___block_739_cmp_zx[20+:1];

_t___block_739_y_sel = _t___block_739_cmp_yx[20+:1]&&~_t___block_739_cmp_zy[20+:1];

_t___block_739_z_sel = _t___block_739_cmp_zx[20+:1]&&_t___block_739_cmp_zy[20+:1];

if (_t___block_739_x_sel) begin
// __block_740
// __block_742
_d___pip_5160_1_40___stage___block_26_v_x = _q___pip_5160_1_40___stage___block_26_v_x+_q___pip_5160_1_40___stage___block_26_s_x;

_d___pip_5160_1_40___block_34_tm_x = _q___pip_5160_1_40___block_34_tm_x+_q___pip_5160_1_40___block_40_dt_x;

// __block_743
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_741
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_744
if (_t___block_739_y_sel) begin
// __block_745
// __block_747
_d___pip_5160_1_40___stage___block_26_v_y = _q___pip_5160_1_40___stage___block_26_v_y+_q___pip_5160_1_40___stage___block_26_s_y;

_d___pip_5160_1_40___block_34_tm_y = _q___pip_5160_1_40___block_34_tm_y+_q___pip_5160_1_40___block_40_dt_y;

// __block_748
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_746
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_749
if (_t___block_739_z_sel) begin
// __block_750
// __block_752
_d___pip_5160_1_40___stage___block_26_v_z = _q___pip_5160_1_40___stage___block_26_v_z+_q___pip_5160_1_40___stage___block_26_s_z;

_d___pip_5160_1_40___block_34_tm_z = _q___pip_5160_1_40___block_34_tm_z+_q___pip_5160_1_40___block_40_dt_z;

// __block_753
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_751
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_754
// end of pipeline stage
_d__full_fsm___pip_5160_1_40 = 1;
_d__idx_fsm___pip_5160_1_40 = _t__stall_fsm___pip_5160_1_40 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_40 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 41
(* full_case *)
case (_q__idx_fsm___pip_5160_1_41)
1: begin
// __stage___block_755
_t___stage___block_755_tex = (_q___pip_5160_1_41___stage___block_26_v_x)^(_q___pip_5160_1_41___stage___block_26_v_y)^(_q___pip_5160_1_41___stage___block_26_v_z);

_t___stage___block_755_vnum0 = {_q___pip_5160_1_41___stage___block_26_v_z[0+:2],_q___pip_5160_1_41___stage___block_26_v_y[0+:2],_q___pip_5160_1_41___stage___block_26_v_x[0+:2]};

_t___stage___block_755_vnum1 = {_q___pip_5160_1_41___stage___block_26_v_z[2+:2],_q___pip_5160_1_41___stage___block_26_v_y[2+:2],_q___pip_5160_1_41___stage___block_26_v_x[2+:2]};

_t___stage___block_755_vnum2 = {_q___pip_5160_1_41___stage___block_26_v_z[4+:2],_q___pip_5160_1_41___stage___block_26_v_y[4+:2],_q___pip_5160_1_41___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_41___stage___block_6_inside&_w_tile[_t___stage___block_755_vnum0+:1]&_w_tile[_t___stage___block_755_vnum1+:1]&_w_tile[_t___stage___block_755_vnum2+:1]) begin
// __block_756
// __block_758
_d___pip_5160_1_41___stage___block_6_clr = _t___stage___block_755_tex;

_d___pip_5160_1_41___stage___block_6_dist = 63;

_d___pip_5160_1_41___stage___block_6_inside = 1;

// __block_759
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_757
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_760
_t___block_760_cmp_yx = _q___pip_5160_1_41___block_34_tm_y-_q___pip_5160_1_41___block_34_tm_x;

_t___block_760_cmp_zx = _q___pip_5160_1_41___block_34_tm_z-_q___pip_5160_1_41___block_34_tm_x;

_t___block_760_cmp_zy = _q___pip_5160_1_41___block_34_tm_z-_q___pip_5160_1_41___block_34_tm_y;

_t___block_760_x_sel = ~_t___block_760_cmp_yx[20+:1]&&~_t___block_760_cmp_zx[20+:1];

_t___block_760_y_sel = _t___block_760_cmp_yx[20+:1]&&~_t___block_760_cmp_zy[20+:1];

_t___block_760_z_sel = _t___block_760_cmp_zx[20+:1]&&_t___block_760_cmp_zy[20+:1];

if (_t___block_760_x_sel) begin
// __block_761
// __block_763
_d___pip_5160_1_41___stage___block_26_v_x = _q___pip_5160_1_41___stage___block_26_v_x+_q___pip_5160_1_41___stage___block_26_s_x;

_d___pip_5160_1_41___block_34_tm_x = _q___pip_5160_1_41___block_34_tm_x+_q___pip_5160_1_41___block_40_dt_x;

// __block_764
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_762
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_765
if (_t___block_760_y_sel) begin
// __block_766
// __block_768
_d___pip_5160_1_41___stage___block_26_v_y = _q___pip_5160_1_41___stage___block_26_v_y+_q___pip_5160_1_41___stage___block_26_s_y;

_d___pip_5160_1_41___block_34_tm_y = _q___pip_5160_1_41___block_34_tm_y+_q___pip_5160_1_41___block_40_dt_y;

// __block_769
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_767
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_770
if (_t___block_760_z_sel) begin
// __block_771
// __block_773
_d___pip_5160_1_41___stage___block_26_v_z = _q___pip_5160_1_41___stage___block_26_v_z+_q___pip_5160_1_41___stage___block_26_s_z;

_d___pip_5160_1_41___block_34_tm_z = _q___pip_5160_1_41___block_34_tm_z+_q___pip_5160_1_41___block_40_dt_z;

// __block_774
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_772
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_775
// end of pipeline stage
_d__full_fsm___pip_5160_1_41 = 1;
_d__idx_fsm___pip_5160_1_41 = _t__stall_fsm___pip_5160_1_41 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_41 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 42
(* full_case *)
case (_q__idx_fsm___pip_5160_1_42)
1: begin
// __stage___block_776
_t___stage___block_776_tex = (_q___pip_5160_1_42___stage___block_26_v_x)^(_q___pip_5160_1_42___stage___block_26_v_y)^(_q___pip_5160_1_42___stage___block_26_v_z);

_t___stage___block_776_vnum0 = {_q___pip_5160_1_42___stage___block_26_v_z[0+:2],_q___pip_5160_1_42___stage___block_26_v_y[0+:2],_q___pip_5160_1_42___stage___block_26_v_x[0+:2]};

_t___stage___block_776_vnum1 = {_q___pip_5160_1_42___stage___block_26_v_z[2+:2],_q___pip_5160_1_42___stage___block_26_v_y[2+:2],_q___pip_5160_1_42___stage___block_26_v_x[2+:2]};

_t___stage___block_776_vnum2 = {_q___pip_5160_1_42___stage___block_26_v_z[4+:2],_q___pip_5160_1_42___stage___block_26_v_y[4+:2],_q___pip_5160_1_42___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_42___stage___block_6_inside&_w_tile[_t___stage___block_776_vnum0+:1]&_w_tile[_t___stage___block_776_vnum1+:1]&_w_tile[_t___stage___block_776_vnum2+:1]) begin
// __block_777
// __block_779
_d___pip_5160_1_42___stage___block_6_clr = _t___stage___block_776_tex;

_d___pip_5160_1_42___stage___block_6_dist = 65;

_d___pip_5160_1_42___stage___block_6_inside = 1;

// __block_780
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_778
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_781
_t___block_781_cmp_yx = _q___pip_5160_1_42___block_34_tm_y-_q___pip_5160_1_42___block_34_tm_x;

_t___block_781_cmp_zx = _q___pip_5160_1_42___block_34_tm_z-_q___pip_5160_1_42___block_34_tm_x;

_t___block_781_cmp_zy = _q___pip_5160_1_42___block_34_tm_z-_q___pip_5160_1_42___block_34_tm_y;

_t___block_781_x_sel = ~_t___block_781_cmp_yx[20+:1]&&~_t___block_781_cmp_zx[20+:1];

_t___block_781_y_sel = _t___block_781_cmp_yx[20+:1]&&~_t___block_781_cmp_zy[20+:1];

_t___block_781_z_sel = _t___block_781_cmp_zx[20+:1]&&_t___block_781_cmp_zy[20+:1];

if (_t___block_781_x_sel) begin
// __block_782
// __block_784
_d___pip_5160_1_42___stage___block_26_v_x = _q___pip_5160_1_42___stage___block_26_v_x+_q___pip_5160_1_42___stage___block_26_s_x;

_d___pip_5160_1_42___block_34_tm_x = _q___pip_5160_1_42___block_34_tm_x+_q___pip_5160_1_42___block_40_dt_x;

// __block_785
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_783
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_786
if (_t___block_781_y_sel) begin
// __block_787
// __block_789
_d___pip_5160_1_42___stage___block_26_v_y = _q___pip_5160_1_42___stage___block_26_v_y+_q___pip_5160_1_42___stage___block_26_s_y;

_d___pip_5160_1_42___block_34_tm_y = _q___pip_5160_1_42___block_34_tm_y+_q___pip_5160_1_42___block_40_dt_y;

// __block_790
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_788
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_791
if (_t___block_781_z_sel) begin
// __block_792
// __block_794
_d___pip_5160_1_42___stage___block_26_v_z = _q___pip_5160_1_42___stage___block_26_v_z+_q___pip_5160_1_42___stage___block_26_s_z;

_d___pip_5160_1_42___block_34_tm_z = _q___pip_5160_1_42___block_34_tm_z+_q___pip_5160_1_42___block_40_dt_z;

// __block_795
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_793
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_796
// end of pipeline stage
_d__full_fsm___pip_5160_1_42 = 1;
_d__idx_fsm___pip_5160_1_42 = _t__stall_fsm___pip_5160_1_42 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_42 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 43
(* full_case *)
case (_q__idx_fsm___pip_5160_1_43)
1: begin
// __stage___block_797
_t___stage___block_797_tex = (_q___pip_5160_1_43___stage___block_26_v_x)^(_q___pip_5160_1_43___stage___block_26_v_y)^(_q___pip_5160_1_43___stage___block_26_v_z);

_t___stage___block_797_vnum0 = {_q___pip_5160_1_43___stage___block_26_v_z[0+:2],_q___pip_5160_1_43___stage___block_26_v_y[0+:2],_q___pip_5160_1_43___stage___block_26_v_x[0+:2]};

_t___stage___block_797_vnum1 = {_q___pip_5160_1_43___stage___block_26_v_z[2+:2],_q___pip_5160_1_43___stage___block_26_v_y[2+:2],_q___pip_5160_1_43___stage___block_26_v_x[2+:2]};

_t___stage___block_797_vnum2 = {_q___pip_5160_1_43___stage___block_26_v_z[4+:2],_q___pip_5160_1_43___stage___block_26_v_y[4+:2],_q___pip_5160_1_43___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_43___stage___block_6_inside&_w_tile[_t___stage___block_797_vnum0+:1]&_w_tile[_t___stage___block_797_vnum1+:1]&_w_tile[_t___stage___block_797_vnum2+:1]) begin
// __block_798
// __block_800
_d___pip_5160_1_43___stage___block_6_clr = _t___stage___block_797_tex;

_d___pip_5160_1_43___stage___block_6_dist = 67;

_d___pip_5160_1_43___stage___block_6_inside = 1;

// __block_801
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_799
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_802
_t___block_802_cmp_yx = _q___pip_5160_1_43___block_34_tm_y-_q___pip_5160_1_43___block_34_tm_x;

_t___block_802_cmp_zx = _q___pip_5160_1_43___block_34_tm_z-_q___pip_5160_1_43___block_34_tm_x;

_t___block_802_cmp_zy = _q___pip_5160_1_43___block_34_tm_z-_q___pip_5160_1_43___block_34_tm_y;

_t___block_802_x_sel = ~_t___block_802_cmp_yx[20+:1]&&~_t___block_802_cmp_zx[20+:1];

_t___block_802_y_sel = _t___block_802_cmp_yx[20+:1]&&~_t___block_802_cmp_zy[20+:1];

_t___block_802_z_sel = _t___block_802_cmp_zx[20+:1]&&_t___block_802_cmp_zy[20+:1];

if (_t___block_802_x_sel) begin
// __block_803
// __block_805
_d___pip_5160_1_43___stage___block_26_v_x = _q___pip_5160_1_43___stage___block_26_v_x+_q___pip_5160_1_43___stage___block_26_s_x;

_d___pip_5160_1_43___block_34_tm_x = _q___pip_5160_1_43___block_34_tm_x+_q___pip_5160_1_43___block_40_dt_x;

// __block_806
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_804
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_807
if (_t___block_802_y_sel) begin
// __block_808
// __block_810
_d___pip_5160_1_43___stage___block_26_v_y = _q___pip_5160_1_43___stage___block_26_v_y+_q___pip_5160_1_43___stage___block_26_s_y;

_d___pip_5160_1_43___block_34_tm_y = _q___pip_5160_1_43___block_34_tm_y+_q___pip_5160_1_43___block_40_dt_y;

// __block_811
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_809
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_812
if (_t___block_802_z_sel) begin
// __block_813
// __block_815
_d___pip_5160_1_43___stage___block_26_v_z = _q___pip_5160_1_43___stage___block_26_v_z+_q___pip_5160_1_43___stage___block_26_s_z;

_d___pip_5160_1_43___block_34_tm_z = _q___pip_5160_1_43___block_34_tm_z+_q___pip_5160_1_43___block_40_dt_z;

// __block_816
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_814
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_817
// end of pipeline stage
_d__full_fsm___pip_5160_1_43 = 1;
_d__idx_fsm___pip_5160_1_43 = _t__stall_fsm___pip_5160_1_43 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_43 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 44
(* full_case *)
case (_q__idx_fsm___pip_5160_1_44)
1: begin
// __stage___block_818
_t___stage___block_818_tex = (_q___pip_5160_1_44___stage___block_26_v_x)^(_q___pip_5160_1_44___stage___block_26_v_y)^(_q___pip_5160_1_44___stage___block_26_v_z);

_t___stage___block_818_vnum0 = {_q___pip_5160_1_44___stage___block_26_v_z[0+:2],_q___pip_5160_1_44___stage___block_26_v_y[0+:2],_q___pip_5160_1_44___stage___block_26_v_x[0+:2]};

_t___stage___block_818_vnum1 = {_q___pip_5160_1_44___stage___block_26_v_z[2+:2],_q___pip_5160_1_44___stage___block_26_v_y[2+:2],_q___pip_5160_1_44___stage___block_26_v_x[2+:2]};

_t___stage___block_818_vnum2 = {_q___pip_5160_1_44___stage___block_26_v_z[4+:2],_q___pip_5160_1_44___stage___block_26_v_y[4+:2],_q___pip_5160_1_44___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_44___stage___block_6_inside&_w_tile[_t___stage___block_818_vnum0+:1]&_w_tile[_t___stage___block_818_vnum1+:1]&_w_tile[_t___stage___block_818_vnum2+:1]) begin
// __block_819
// __block_821
_d___pip_5160_1_44___stage___block_6_clr = _t___stage___block_818_tex;

_d___pip_5160_1_44___stage___block_6_dist = 69;

_d___pip_5160_1_44___stage___block_6_inside = 1;

// __block_822
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_820
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_823
_t___block_823_cmp_yx = _q___pip_5160_1_44___block_34_tm_y-_q___pip_5160_1_44___block_34_tm_x;

_t___block_823_cmp_zx = _q___pip_5160_1_44___block_34_tm_z-_q___pip_5160_1_44___block_34_tm_x;

_t___block_823_cmp_zy = _q___pip_5160_1_44___block_34_tm_z-_q___pip_5160_1_44___block_34_tm_y;

_t___block_823_x_sel = ~_t___block_823_cmp_yx[20+:1]&&~_t___block_823_cmp_zx[20+:1];

_t___block_823_y_sel = _t___block_823_cmp_yx[20+:1]&&~_t___block_823_cmp_zy[20+:1];

_t___block_823_z_sel = _t___block_823_cmp_zx[20+:1]&&_t___block_823_cmp_zy[20+:1];

if (_t___block_823_x_sel) begin
// __block_824
// __block_826
_d___pip_5160_1_44___stage___block_26_v_x = _q___pip_5160_1_44___stage___block_26_v_x+_q___pip_5160_1_44___stage___block_26_s_x;

_d___pip_5160_1_44___block_34_tm_x = _q___pip_5160_1_44___block_34_tm_x+_q___pip_5160_1_44___block_40_dt_x;

// __block_827
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_825
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_828
if (_t___block_823_y_sel) begin
// __block_829
// __block_831
_d___pip_5160_1_44___stage___block_26_v_y = _q___pip_5160_1_44___stage___block_26_v_y+_q___pip_5160_1_44___stage___block_26_s_y;

_d___pip_5160_1_44___block_34_tm_y = _q___pip_5160_1_44___block_34_tm_y+_q___pip_5160_1_44___block_40_dt_y;

// __block_832
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_830
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_833
if (_t___block_823_z_sel) begin
// __block_834
// __block_836
_d___pip_5160_1_44___stage___block_26_v_z = _q___pip_5160_1_44___stage___block_26_v_z+_q___pip_5160_1_44___stage___block_26_s_z;

_d___pip_5160_1_44___block_34_tm_z = _q___pip_5160_1_44___block_34_tm_z+_q___pip_5160_1_44___block_40_dt_z;

// __block_837
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_835
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_838
// end of pipeline stage
_d__full_fsm___pip_5160_1_44 = 1;
_d__idx_fsm___pip_5160_1_44 = _t__stall_fsm___pip_5160_1_44 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_44 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 45
(* full_case *)
case (_q__idx_fsm___pip_5160_1_45)
1: begin
// __stage___block_839
_t___stage___block_839_tex = (_q___pip_5160_1_45___stage___block_26_v_x)^(_q___pip_5160_1_45___stage___block_26_v_y)^(_q___pip_5160_1_45___stage___block_26_v_z);

_t___stage___block_839_vnum0 = {_q___pip_5160_1_45___stage___block_26_v_z[0+:2],_q___pip_5160_1_45___stage___block_26_v_y[0+:2],_q___pip_5160_1_45___stage___block_26_v_x[0+:2]};

_t___stage___block_839_vnum1 = {_q___pip_5160_1_45___stage___block_26_v_z[2+:2],_q___pip_5160_1_45___stage___block_26_v_y[2+:2],_q___pip_5160_1_45___stage___block_26_v_x[2+:2]};

_t___stage___block_839_vnum2 = {_q___pip_5160_1_45___stage___block_26_v_z[4+:2],_q___pip_5160_1_45___stage___block_26_v_y[4+:2],_q___pip_5160_1_45___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_45___stage___block_6_inside&_w_tile[_t___stage___block_839_vnum0+:1]&_w_tile[_t___stage___block_839_vnum1+:1]&_w_tile[_t___stage___block_839_vnum2+:1]) begin
// __block_840
// __block_842
_d___pip_5160_1_45___stage___block_6_clr = _t___stage___block_839_tex;

_d___pip_5160_1_45___stage___block_6_dist = 70;

_d___pip_5160_1_45___stage___block_6_inside = 1;

// __block_843
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_841
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_844
_t___block_844_cmp_yx = _q___pip_5160_1_45___block_34_tm_y-_q___pip_5160_1_45___block_34_tm_x;

_t___block_844_cmp_zx = _q___pip_5160_1_45___block_34_tm_z-_q___pip_5160_1_45___block_34_tm_x;

_t___block_844_cmp_zy = _q___pip_5160_1_45___block_34_tm_z-_q___pip_5160_1_45___block_34_tm_y;

_t___block_844_x_sel = ~_t___block_844_cmp_yx[20+:1]&&~_t___block_844_cmp_zx[20+:1];

_t___block_844_y_sel = _t___block_844_cmp_yx[20+:1]&&~_t___block_844_cmp_zy[20+:1];

_t___block_844_z_sel = _t___block_844_cmp_zx[20+:1]&&_t___block_844_cmp_zy[20+:1];

if (_t___block_844_x_sel) begin
// __block_845
// __block_847
_d___pip_5160_1_45___stage___block_26_v_x = _q___pip_5160_1_45___stage___block_26_v_x+_q___pip_5160_1_45___stage___block_26_s_x;

_d___pip_5160_1_45___block_34_tm_x = _q___pip_5160_1_45___block_34_tm_x+_q___pip_5160_1_45___block_40_dt_x;

// __block_848
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_846
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_849
if (_t___block_844_y_sel) begin
// __block_850
// __block_852
_d___pip_5160_1_45___stage___block_26_v_y = _q___pip_5160_1_45___stage___block_26_v_y+_q___pip_5160_1_45___stage___block_26_s_y;

_d___pip_5160_1_45___block_34_tm_y = _q___pip_5160_1_45___block_34_tm_y+_q___pip_5160_1_45___block_40_dt_y;

// __block_853
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_851
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_854
if (_t___block_844_z_sel) begin
// __block_855
// __block_857
_d___pip_5160_1_45___stage___block_26_v_z = _q___pip_5160_1_45___stage___block_26_v_z+_q___pip_5160_1_45___stage___block_26_s_z;

_d___pip_5160_1_45___block_34_tm_z = _q___pip_5160_1_45___block_34_tm_z+_q___pip_5160_1_45___block_40_dt_z;

// __block_858
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_856
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_859
// end of pipeline stage
_d__full_fsm___pip_5160_1_45 = 1;
_d__idx_fsm___pip_5160_1_45 = _t__stall_fsm___pip_5160_1_45 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_45 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 46
(* full_case *)
case (_q__idx_fsm___pip_5160_1_46)
1: begin
// __stage___block_860
_t___stage___block_860_tex = (_q___pip_5160_1_46___stage___block_26_v_x)^(_q___pip_5160_1_46___stage___block_26_v_y)^(_q___pip_5160_1_46___stage___block_26_v_z);

_t___stage___block_860_vnum0 = {_q___pip_5160_1_46___stage___block_26_v_z[0+:2],_q___pip_5160_1_46___stage___block_26_v_y[0+:2],_q___pip_5160_1_46___stage___block_26_v_x[0+:2]};

_t___stage___block_860_vnum1 = {_q___pip_5160_1_46___stage___block_26_v_z[2+:2],_q___pip_5160_1_46___stage___block_26_v_y[2+:2],_q___pip_5160_1_46___stage___block_26_v_x[2+:2]};

_t___stage___block_860_vnum2 = {_q___pip_5160_1_46___stage___block_26_v_z[4+:2],_q___pip_5160_1_46___stage___block_26_v_y[4+:2],_q___pip_5160_1_46___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_46___stage___block_6_inside&_w_tile[_t___stage___block_860_vnum0+:1]&_w_tile[_t___stage___block_860_vnum1+:1]&_w_tile[_t___stage___block_860_vnum2+:1]) begin
// __block_861
// __block_863
_d___pip_5160_1_46___stage___block_6_clr = _t___stage___block_860_tex;

_d___pip_5160_1_46___stage___block_6_dist = 72;

_d___pip_5160_1_46___stage___block_6_inside = 1;

// __block_864
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_862
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_865
_t___block_865_cmp_yx = _q___pip_5160_1_46___block_34_tm_y-_q___pip_5160_1_46___block_34_tm_x;

_t___block_865_cmp_zx = _q___pip_5160_1_46___block_34_tm_z-_q___pip_5160_1_46___block_34_tm_x;

_t___block_865_cmp_zy = _q___pip_5160_1_46___block_34_tm_z-_q___pip_5160_1_46___block_34_tm_y;

_t___block_865_x_sel = ~_t___block_865_cmp_yx[20+:1]&&~_t___block_865_cmp_zx[20+:1];

_t___block_865_y_sel = _t___block_865_cmp_yx[20+:1]&&~_t___block_865_cmp_zy[20+:1];

_t___block_865_z_sel = _t___block_865_cmp_zx[20+:1]&&_t___block_865_cmp_zy[20+:1];

if (_t___block_865_x_sel) begin
// __block_866
// __block_868
_d___pip_5160_1_46___stage___block_26_v_x = _q___pip_5160_1_46___stage___block_26_v_x+_q___pip_5160_1_46___stage___block_26_s_x;

_d___pip_5160_1_46___block_34_tm_x = _q___pip_5160_1_46___block_34_tm_x+_q___pip_5160_1_46___block_40_dt_x;

// __block_869
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_867
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_870
if (_t___block_865_y_sel) begin
// __block_871
// __block_873
_d___pip_5160_1_46___stage___block_26_v_y = _q___pip_5160_1_46___stage___block_26_v_y+_q___pip_5160_1_46___stage___block_26_s_y;

_d___pip_5160_1_46___block_34_tm_y = _q___pip_5160_1_46___block_34_tm_y+_q___pip_5160_1_46___block_40_dt_y;

// __block_874
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_872
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_875
if (_t___block_865_z_sel) begin
// __block_876
// __block_878
_d___pip_5160_1_46___stage___block_26_v_z = _q___pip_5160_1_46___stage___block_26_v_z+_q___pip_5160_1_46___stage___block_26_s_z;

_d___pip_5160_1_46___block_34_tm_z = _q___pip_5160_1_46___block_34_tm_z+_q___pip_5160_1_46___block_40_dt_z;

// __block_879
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_877
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_880
// end of pipeline stage
_d__full_fsm___pip_5160_1_46 = 1;
_d__idx_fsm___pip_5160_1_46 = _t__stall_fsm___pip_5160_1_46 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_46 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 47
(* full_case *)
case (_q__idx_fsm___pip_5160_1_47)
1: begin
// __stage___block_881
_t___stage___block_881_tex = (_q___pip_5160_1_47___stage___block_26_v_x)^(_q___pip_5160_1_47___stage___block_26_v_y)^(_q___pip_5160_1_47___stage___block_26_v_z);

_t___stage___block_881_vnum0 = {_q___pip_5160_1_47___stage___block_26_v_z[0+:2],_q___pip_5160_1_47___stage___block_26_v_y[0+:2],_q___pip_5160_1_47___stage___block_26_v_x[0+:2]};

_t___stage___block_881_vnum1 = {_q___pip_5160_1_47___stage___block_26_v_z[2+:2],_q___pip_5160_1_47___stage___block_26_v_y[2+:2],_q___pip_5160_1_47___stage___block_26_v_x[2+:2]};

_t___stage___block_881_vnum2 = {_q___pip_5160_1_47___stage___block_26_v_z[4+:2],_q___pip_5160_1_47___stage___block_26_v_y[4+:2],_q___pip_5160_1_47___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_47___stage___block_6_inside&_w_tile[_t___stage___block_881_vnum0+:1]&_w_tile[_t___stage___block_881_vnum1+:1]&_w_tile[_t___stage___block_881_vnum2+:1]) begin
// __block_882
// __block_884
_d___pip_5160_1_47___stage___block_6_clr = _t___stage___block_881_tex;

_d___pip_5160_1_47___stage___block_6_dist = 74;

_d___pip_5160_1_47___stage___block_6_inside = 1;

// __block_885
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_883
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_886
_t___block_886_cmp_yx = _q___pip_5160_1_47___block_34_tm_y-_q___pip_5160_1_47___block_34_tm_x;

_t___block_886_cmp_zx = _q___pip_5160_1_47___block_34_tm_z-_q___pip_5160_1_47___block_34_tm_x;

_t___block_886_cmp_zy = _q___pip_5160_1_47___block_34_tm_z-_q___pip_5160_1_47___block_34_tm_y;

_t___block_886_x_sel = ~_t___block_886_cmp_yx[20+:1]&&~_t___block_886_cmp_zx[20+:1];

_t___block_886_y_sel = _t___block_886_cmp_yx[20+:1]&&~_t___block_886_cmp_zy[20+:1];

_t___block_886_z_sel = _t___block_886_cmp_zx[20+:1]&&_t___block_886_cmp_zy[20+:1];

if (_t___block_886_x_sel) begin
// __block_887
// __block_889
_d___pip_5160_1_47___stage___block_26_v_x = _q___pip_5160_1_47___stage___block_26_v_x+_q___pip_5160_1_47___stage___block_26_s_x;

_d___pip_5160_1_47___block_34_tm_x = _q___pip_5160_1_47___block_34_tm_x+_q___pip_5160_1_47___block_40_dt_x;

// __block_890
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_888
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_891
if (_t___block_886_y_sel) begin
// __block_892
// __block_894
_d___pip_5160_1_47___stage___block_26_v_y = _q___pip_5160_1_47___stage___block_26_v_y+_q___pip_5160_1_47___stage___block_26_s_y;

_d___pip_5160_1_47___block_34_tm_y = _q___pip_5160_1_47___block_34_tm_y+_q___pip_5160_1_47___block_40_dt_y;

// __block_895
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_893
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_896
if (_t___block_886_z_sel) begin
// __block_897
// __block_899
_d___pip_5160_1_47___stage___block_26_v_z = _q___pip_5160_1_47___stage___block_26_v_z+_q___pip_5160_1_47___stage___block_26_s_z;

_d___pip_5160_1_47___block_34_tm_z = _q___pip_5160_1_47___block_34_tm_z+_q___pip_5160_1_47___block_40_dt_z;

// __block_900
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_898
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_901
// end of pipeline stage
_d__full_fsm___pip_5160_1_47 = 1;
_d__idx_fsm___pip_5160_1_47 = _t__stall_fsm___pip_5160_1_47 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_47 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 48
(* full_case *)
case (_q__idx_fsm___pip_5160_1_48)
1: begin
// __stage___block_902
_t___stage___block_902_tex = (_q___pip_5160_1_48___stage___block_26_v_x)^(_q___pip_5160_1_48___stage___block_26_v_y)^(_q___pip_5160_1_48___stage___block_26_v_z);

_t___stage___block_902_vnum0 = {_q___pip_5160_1_48___stage___block_26_v_z[0+:2],_q___pip_5160_1_48___stage___block_26_v_y[0+:2],_q___pip_5160_1_48___stage___block_26_v_x[0+:2]};

_t___stage___block_902_vnum1 = {_q___pip_5160_1_48___stage___block_26_v_z[2+:2],_q___pip_5160_1_48___stage___block_26_v_y[2+:2],_q___pip_5160_1_48___stage___block_26_v_x[2+:2]};

_t___stage___block_902_vnum2 = {_q___pip_5160_1_48___stage___block_26_v_z[4+:2],_q___pip_5160_1_48___stage___block_26_v_y[4+:2],_q___pip_5160_1_48___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_48___stage___block_6_inside&_w_tile[_t___stage___block_902_vnum0+:1]&_w_tile[_t___stage___block_902_vnum1+:1]&_w_tile[_t___stage___block_902_vnum2+:1]) begin
// __block_903
// __block_905
_d___pip_5160_1_48___stage___block_6_clr = _t___stage___block_902_tex;

_d___pip_5160_1_48___stage___block_6_dist = 76;

_d___pip_5160_1_48___stage___block_6_inside = 1;

// __block_906
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_904
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_907
_t___block_907_cmp_yx = _q___pip_5160_1_48___block_34_tm_y-_q___pip_5160_1_48___block_34_tm_x;

_t___block_907_cmp_zx = _q___pip_5160_1_48___block_34_tm_z-_q___pip_5160_1_48___block_34_tm_x;

_t___block_907_cmp_zy = _q___pip_5160_1_48___block_34_tm_z-_q___pip_5160_1_48___block_34_tm_y;

_t___block_907_x_sel = ~_t___block_907_cmp_yx[20+:1]&&~_t___block_907_cmp_zx[20+:1];

_t___block_907_y_sel = _t___block_907_cmp_yx[20+:1]&&~_t___block_907_cmp_zy[20+:1];

_t___block_907_z_sel = _t___block_907_cmp_zx[20+:1]&&_t___block_907_cmp_zy[20+:1];

if (_t___block_907_x_sel) begin
// __block_908
// __block_910
_d___pip_5160_1_48___stage___block_26_v_x = _q___pip_5160_1_48___stage___block_26_v_x+_q___pip_5160_1_48___stage___block_26_s_x;

_d___pip_5160_1_48___block_34_tm_x = _q___pip_5160_1_48___block_34_tm_x+_q___pip_5160_1_48___block_40_dt_x;

// __block_911
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_909
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_912
if (_t___block_907_y_sel) begin
// __block_913
// __block_915
_d___pip_5160_1_48___stage___block_26_v_y = _q___pip_5160_1_48___stage___block_26_v_y+_q___pip_5160_1_48___stage___block_26_s_y;

_d___pip_5160_1_48___block_34_tm_y = _q___pip_5160_1_48___block_34_tm_y+_q___pip_5160_1_48___block_40_dt_y;

// __block_916
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_914
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_917
if (_t___block_907_z_sel) begin
// __block_918
// __block_920
_d___pip_5160_1_48___stage___block_26_v_z = _q___pip_5160_1_48___stage___block_26_v_z+_q___pip_5160_1_48___stage___block_26_s_z;

_d___pip_5160_1_48___block_34_tm_z = _q___pip_5160_1_48___block_34_tm_z+_q___pip_5160_1_48___block_40_dt_z;

// __block_921
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_919
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_922
// end of pipeline stage
_d__full_fsm___pip_5160_1_48 = 1;
_d__idx_fsm___pip_5160_1_48 = _t__stall_fsm___pip_5160_1_48 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_48 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 49
(* full_case *)
case (_q__idx_fsm___pip_5160_1_49)
1: begin
// __stage___block_923
_t___stage___block_923_tex = (_q___pip_5160_1_49___stage___block_26_v_x)^(_q___pip_5160_1_49___stage___block_26_v_y)^(_q___pip_5160_1_49___stage___block_26_v_z);

_t___stage___block_923_vnum0 = {_q___pip_5160_1_49___stage___block_26_v_z[0+:2],_q___pip_5160_1_49___stage___block_26_v_y[0+:2],_q___pip_5160_1_49___stage___block_26_v_x[0+:2]};

_t___stage___block_923_vnum1 = {_q___pip_5160_1_49___stage___block_26_v_z[2+:2],_q___pip_5160_1_49___stage___block_26_v_y[2+:2],_q___pip_5160_1_49___stage___block_26_v_x[2+:2]};

_t___stage___block_923_vnum2 = {_q___pip_5160_1_49___stage___block_26_v_z[4+:2],_q___pip_5160_1_49___stage___block_26_v_y[4+:2],_q___pip_5160_1_49___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_49___stage___block_6_inside&_w_tile[_t___stage___block_923_vnum0+:1]&_w_tile[_t___stage___block_923_vnum1+:1]&_w_tile[_t___stage___block_923_vnum2+:1]) begin
// __block_924
// __block_926
_d___pip_5160_1_49___stage___block_6_clr = _t___stage___block_923_tex;

_d___pip_5160_1_49___stage___block_6_dist = 78;

_d___pip_5160_1_49___stage___block_6_inside = 1;

// __block_927
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_925
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_928
_t___block_928_cmp_yx = _q___pip_5160_1_49___block_34_tm_y-_q___pip_5160_1_49___block_34_tm_x;

_t___block_928_cmp_zx = _q___pip_5160_1_49___block_34_tm_z-_q___pip_5160_1_49___block_34_tm_x;

_t___block_928_cmp_zy = _q___pip_5160_1_49___block_34_tm_z-_q___pip_5160_1_49___block_34_tm_y;

_t___block_928_x_sel = ~_t___block_928_cmp_yx[20+:1]&&~_t___block_928_cmp_zx[20+:1];

_t___block_928_y_sel = _t___block_928_cmp_yx[20+:1]&&~_t___block_928_cmp_zy[20+:1];

_t___block_928_z_sel = _t___block_928_cmp_zx[20+:1]&&_t___block_928_cmp_zy[20+:1];

if (_t___block_928_x_sel) begin
// __block_929
// __block_931
_d___pip_5160_1_49___stage___block_26_v_x = _q___pip_5160_1_49___stage___block_26_v_x+_q___pip_5160_1_49___stage___block_26_s_x;

_d___pip_5160_1_49___block_34_tm_x = _q___pip_5160_1_49___block_34_tm_x+_q___pip_5160_1_49___block_40_dt_x;

// __block_932
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_930
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_933
if (_t___block_928_y_sel) begin
// __block_934
// __block_936
_d___pip_5160_1_49___stage___block_26_v_y = _q___pip_5160_1_49___stage___block_26_v_y+_q___pip_5160_1_49___stage___block_26_s_y;

_d___pip_5160_1_49___block_34_tm_y = _q___pip_5160_1_49___block_34_tm_y+_q___pip_5160_1_49___block_40_dt_y;

// __block_937
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_935
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_938
if (_t___block_928_z_sel) begin
// __block_939
// __block_941
_d___pip_5160_1_49___stage___block_26_v_z = _q___pip_5160_1_49___stage___block_26_v_z+_q___pip_5160_1_49___stage___block_26_s_z;

_d___pip_5160_1_49___block_34_tm_z = _q___pip_5160_1_49___block_34_tm_z+_q___pip_5160_1_49___block_40_dt_z;

// __block_942
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_940
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_943
// end of pipeline stage
_d__full_fsm___pip_5160_1_49 = 1;
_d__idx_fsm___pip_5160_1_49 = _t__stall_fsm___pip_5160_1_49 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_49 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 50
(* full_case *)
case (_q__idx_fsm___pip_5160_1_50)
1: begin
// __stage___block_944
_t___stage___block_944_tex = (_q___pip_5160_1_50___stage___block_26_v_x)^(_q___pip_5160_1_50___stage___block_26_v_y)^(_q___pip_5160_1_50___stage___block_26_v_z);

_t___stage___block_944_vnum0 = {_q___pip_5160_1_50___stage___block_26_v_z[0+:2],_q___pip_5160_1_50___stage___block_26_v_y[0+:2],_q___pip_5160_1_50___stage___block_26_v_x[0+:2]};

_t___stage___block_944_vnum1 = {_q___pip_5160_1_50___stage___block_26_v_z[2+:2],_q___pip_5160_1_50___stage___block_26_v_y[2+:2],_q___pip_5160_1_50___stage___block_26_v_x[2+:2]};

_t___stage___block_944_vnum2 = {_q___pip_5160_1_50___stage___block_26_v_z[4+:2],_q___pip_5160_1_50___stage___block_26_v_y[4+:2],_q___pip_5160_1_50___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_50___stage___block_6_inside&_w_tile[_t___stage___block_944_vnum0+:1]&_w_tile[_t___stage___block_944_vnum1+:1]&_w_tile[_t___stage___block_944_vnum2+:1]) begin
// __block_945
// __block_947
_d___pip_5160_1_50___stage___block_6_clr = _t___stage___block_944_tex;

_d___pip_5160_1_50___stage___block_6_dist = 80;

_d___pip_5160_1_50___stage___block_6_inside = 1;

// __block_948
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_946
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_949
_t___block_949_cmp_yx = _q___pip_5160_1_50___block_34_tm_y-_q___pip_5160_1_50___block_34_tm_x;

_t___block_949_cmp_zx = _q___pip_5160_1_50___block_34_tm_z-_q___pip_5160_1_50___block_34_tm_x;

_t___block_949_cmp_zy = _q___pip_5160_1_50___block_34_tm_z-_q___pip_5160_1_50___block_34_tm_y;

_t___block_949_x_sel = ~_t___block_949_cmp_yx[20+:1]&&~_t___block_949_cmp_zx[20+:1];

_t___block_949_y_sel = _t___block_949_cmp_yx[20+:1]&&~_t___block_949_cmp_zy[20+:1];

_t___block_949_z_sel = _t___block_949_cmp_zx[20+:1]&&_t___block_949_cmp_zy[20+:1];

if (_t___block_949_x_sel) begin
// __block_950
// __block_952
_d___pip_5160_1_50___stage___block_26_v_x = _q___pip_5160_1_50___stage___block_26_v_x+_q___pip_5160_1_50___stage___block_26_s_x;

_d___pip_5160_1_50___block_34_tm_x = _q___pip_5160_1_50___block_34_tm_x+_q___pip_5160_1_50___block_40_dt_x;

// __block_953
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_951
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_954
if (_t___block_949_y_sel) begin
// __block_955
// __block_957
_d___pip_5160_1_50___stage___block_26_v_y = _q___pip_5160_1_50___stage___block_26_v_y+_q___pip_5160_1_50___stage___block_26_s_y;

_d___pip_5160_1_50___block_34_tm_y = _q___pip_5160_1_50___block_34_tm_y+_q___pip_5160_1_50___block_40_dt_y;

// __block_958
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_956
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_959
if (_t___block_949_z_sel) begin
// __block_960
// __block_962
_d___pip_5160_1_50___stage___block_26_v_z = _q___pip_5160_1_50___stage___block_26_v_z+_q___pip_5160_1_50___stage___block_26_s_z;

_d___pip_5160_1_50___block_34_tm_z = _q___pip_5160_1_50___block_34_tm_z+_q___pip_5160_1_50___block_40_dt_z;

// __block_963
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_961
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_964
// end of pipeline stage
_d__full_fsm___pip_5160_1_50 = 1;
_d__idx_fsm___pip_5160_1_50 = _t__stall_fsm___pip_5160_1_50 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_50 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 51
(* full_case *)
case (_q__idx_fsm___pip_5160_1_51)
1: begin
// __stage___block_965
_t___stage___block_965_tex = (_q___pip_5160_1_51___stage___block_26_v_x)^(_q___pip_5160_1_51___stage___block_26_v_y)^(_q___pip_5160_1_51___stage___block_26_v_z);

_t___stage___block_965_vnum0 = {_q___pip_5160_1_51___stage___block_26_v_z[0+:2],_q___pip_5160_1_51___stage___block_26_v_y[0+:2],_q___pip_5160_1_51___stage___block_26_v_x[0+:2]};

_t___stage___block_965_vnum1 = {_q___pip_5160_1_51___stage___block_26_v_z[2+:2],_q___pip_5160_1_51___stage___block_26_v_y[2+:2],_q___pip_5160_1_51___stage___block_26_v_x[2+:2]};

_t___stage___block_965_vnum2 = {_q___pip_5160_1_51___stage___block_26_v_z[4+:2],_q___pip_5160_1_51___stage___block_26_v_y[4+:2],_q___pip_5160_1_51___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_51___stage___block_6_inside&_w_tile[_t___stage___block_965_vnum0+:1]&_w_tile[_t___stage___block_965_vnum1+:1]&_w_tile[_t___stage___block_965_vnum2+:1]) begin
// __block_966
// __block_968
_d___pip_5160_1_51___stage___block_6_clr = _t___stage___block_965_tex;

_d___pip_5160_1_51___stage___block_6_dist = 82;

_d___pip_5160_1_51___stage___block_6_inside = 1;

// __block_969
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_967
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_970
_t___block_970_cmp_yx = _q___pip_5160_1_51___block_34_tm_y-_q___pip_5160_1_51___block_34_tm_x;

_t___block_970_cmp_zx = _q___pip_5160_1_51___block_34_tm_z-_q___pip_5160_1_51___block_34_tm_x;

_t___block_970_cmp_zy = _q___pip_5160_1_51___block_34_tm_z-_q___pip_5160_1_51___block_34_tm_y;

_t___block_970_x_sel = ~_t___block_970_cmp_yx[20+:1]&&~_t___block_970_cmp_zx[20+:1];

_t___block_970_y_sel = _t___block_970_cmp_yx[20+:1]&&~_t___block_970_cmp_zy[20+:1];

_t___block_970_z_sel = _t___block_970_cmp_zx[20+:1]&&_t___block_970_cmp_zy[20+:1];

if (_t___block_970_x_sel) begin
// __block_971
// __block_973
_d___pip_5160_1_51___stage___block_26_v_x = _q___pip_5160_1_51___stage___block_26_v_x+_q___pip_5160_1_51___stage___block_26_s_x;

_d___pip_5160_1_51___block_34_tm_x = _q___pip_5160_1_51___block_34_tm_x+_q___pip_5160_1_51___block_40_dt_x;

// __block_974
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_972
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_975
if (_t___block_970_y_sel) begin
// __block_976
// __block_978
_d___pip_5160_1_51___stage___block_26_v_y = _q___pip_5160_1_51___stage___block_26_v_y+_q___pip_5160_1_51___stage___block_26_s_y;

_d___pip_5160_1_51___block_34_tm_y = _q___pip_5160_1_51___block_34_tm_y+_q___pip_5160_1_51___block_40_dt_y;

// __block_979
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_977
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_980
if (_t___block_970_z_sel) begin
// __block_981
// __block_983
_d___pip_5160_1_51___stage___block_26_v_z = _q___pip_5160_1_51___stage___block_26_v_z+_q___pip_5160_1_51___stage___block_26_s_z;

_d___pip_5160_1_51___block_34_tm_z = _q___pip_5160_1_51___block_34_tm_z+_q___pip_5160_1_51___block_40_dt_z;

// __block_984
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_982
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_985
// end of pipeline stage
_d__full_fsm___pip_5160_1_51 = 1;
_d__idx_fsm___pip_5160_1_51 = _t__stall_fsm___pip_5160_1_51 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_51 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 52
(* full_case *)
case (_q__idx_fsm___pip_5160_1_52)
1: begin
// __stage___block_986
_t___stage___block_986_tex = (_q___pip_5160_1_52___stage___block_26_v_x)^(_q___pip_5160_1_52___stage___block_26_v_y)^(_q___pip_5160_1_52___stage___block_26_v_z);

_t___stage___block_986_vnum0 = {_q___pip_5160_1_52___stage___block_26_v_z[0+:2],_q___pip_5160_1_52___stage___block_26_v_y[0+:2],_q___pip_5160_1_52___stage___block_26_v_x[0+:2]};

_t___stage___block_986_vnum1 = {_q___pip_5160_1_52___stage___block_26_v_z[2+:2],_q___pip_5160_1_52___stage___block_26_v_y[2+:2],_q___pip_5160_1_52___stage___block_26_v_x[2+:2]};

_t___stage___block_986_vnum2 = {_q___pip_5160_1_52___stage___block_26_v_z[4+:2],_q___pip_5160_1_52___stage___block_26_v_y[4+:2],_q___pip_5160_1_52___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_52___stage___block_6_inside&_w_tile[_t___stage___block_986_vnum0+:1]&_w_tile[_t___stage___block_986_vnum1+:1]&_w_tile[_t___stage___block_986_vnum2+:1]) begin
// __block_987
// __block_989
_d___pip_5160_1_52___stage___block_6_clr = _t___stage___block_986_tex;

_d___pip_5160_1_52___stage___block_6_dist = 84;

_d___pip_5160_1_52___stage___block_6_inside = 1;

// __block_990
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_988
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_991
_t___block_991_cmp_yx = _q___pip_5160_1_52___block_34_tm_y-_q___pip_5160_1_52___block_34_tm_x;

_t___block_991_cmp_zx = _q___pip_5160_1_52___block_34_tm_z-_q___pip_5160_1_52___block_34_tm_x;

_t___block_991_cmp_zy = _q___pip_5160_1_52___block_34_tm_z-_q___pip_5160_1_52___block_34_tm_y;

_t___block_991_x_sel = ~_t___block_991_cmp_yx[20+:1]&&~_t___block_991_cmp_zx[20+:1];

_t___block_991_y_sel = _t___block_991_cmp_yx[20+:1]&&~_t___block_991_cmp_zy[20+:1];

_t___block_991_z_sel = _t___block_991_cmp_zx[20+:1]&&_t___block_991_cmp_zy[20+:1];

if (_t___block_991_x_sel) begin
// __block_992
// __block_994
_d___pip_5160_1_52___stage___block_26_v_x = _q___pip_5160_1_52___stage___block_26_v_x+_q___pip_5160_1_52___stage___block_26_s_x;

_d___pip_5160_1_52___block_34_tm_x = _q___pip_5160_1_52___block_34_tm_x+_q___pip_5160_1_52___block_40_dt_x;

// __block_995
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_993
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_996
if (_t___block_991_y_sel) begin
// __block_997
// __block_999
_d___pip_5160_1_52___stage___block_26_v_y = _q___pip_5160_1_52___stage___block_26_v_y+_q___pip_5160_1_52___stage___block_26_s_y;

_d___pip_5160_1_52___block_34_tm_y = _q___pip_5160_1_52___block_34_tm_y+_q___pip_5160_1_52___block_40_dt_y;

// __block_1000
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_998
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1001
if (_t___block_991_z_sel) begin
// __block_1002
// __block_1004
_d___pip_5160_1_52___stage___block_26_v_z = _q___pip_5160_1_52___stage___block_26_v_z+_q___pip_5160_1_52___stage___block_26_s_z;

_d___pip_5160_1_52___block_34_tm_z = _q___pip_5160_1_52___block_34_tm_z+_q___pip_5160_1_52___block_40_dt_z;

// __block_1005
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1003
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1006
// end of pipeline stage
_d__full_fsm___pip_5160_1_52 = 1;
_d__idx_fsm___pip_5160_1_52 = _t__stall_fsm___pip_5160_1_52 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_52 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 53
(* full_case *)
case (_q__idx_fsm___pip_5160_1_53)
1: begin
// __stage___block_1007
_t___stage___block_1007_tex = (_q___pip_5160_1_53___stage___block_26_v_x)^(_q___pip_5160_1_53___stage___block_26_v_y)^(_q___pip_5160_1_53___stage___block_26_v_z);

_t___stage___block_1007_vnum0 = {_q___pip_5160_1_53___stage___block_26_v_z[0+:2],_q___pip_5160_1_53___stage___block_26_v_y[0+:2],_q___pip_5160_1_53___stage___block_26_v_x[0+:2]};

_t___stage___block_1007_vnum1 = {_q___pip_5160_1_53___stage___block_26_v_z[2+:2],_q___pip_5160_1_53___stage___block_26_v_y[2+:2],_q___pip_5160_1_53___stage___block_26_v_x[2+:2]};

_t___stage___block_1007_vnum2 = {_q___pip_5160_1_53___stage___block_26_v_z[4+:2],_q___pip_5160_1_53___stage___block_26_v_y[4+:2],_q___pip_5160_1_53___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_53___stage___block_6_inside&_w_tile[_t___stage___block_1007_vnum0+:1]&_w_tile[_t___stage___block_1007_vnum1+:1]&_w_tile[_t___stage___block_1007_vnum2+:1]) begin
// __block_1008
// __block_1010
_d___pip_5160_1_53___stage___block_6_clr = _t___stage___block_1007_tex;

_d___pip_5160_1_53___stage___block_6_dist = 85;

_d___pip_5160_1_53___stage___block_6_inside = 1;

// __block_1011
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1009
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1012
_t___block_1012_cmp_yx = _q___pip_5160_1_53___block_34_tm_y-_q___pip_5160_1_53___block_34_tm_x;

_t___block_1012_cmp_zx = _q___pip_5160_1_53___block_34_tm_z-_q___pip_5160_1_53___block_34_tm_x;

_t___block_1012_cmp_zy = _q___pip_5160_1_53___block_34_tm_z-_q___pip_5160_1_53___block_34_tm_y;

_t___block_1012_x_sel = ~_t___block_1012_cmp_yx[20+:1]&&~_t___block_1012_cmp_zx[20+:1];

_t___block_1012_y_sel = _t___block_1012_cmp_yx[20+:1]&&~_t___block_1012_cmp_zy[20+:1];

_t___block_1012_z_sel = _t___block_1012_cmp_zx[20+:1]&&_t___block_1012_cmp_zy[20+:1];

if (_t___block_1012_x_sel) begin
// __block_1013
// __block_1015
_d___pip_5160_1_53___stage___block_26_v_x = _q___pip_5160_1_53___stage___block_26_v_x+_q___pip_5160_1_53___stage___block_26_s_x;

_d___pip_5160_1_53___block_34_tm_x = _q___pip_5160_1_53___block_34_tm_x+_q___pip_5160_1_53___block_40_dt_x;

// __block_1016
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1014
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1017
if (_t___block_1012_y_sel) begin
// __block_1018
// __block_1020
_d___pip_5160_1_53___stage___block_26_v_y = _q___pip_5160_1_53___stage___block_26_v_y+_q___pip_5160_1_53___stage___block_26_s_y;

_d___pip_5160_1_53___block_34_tm_y = _q___pip_5160_1_53___block_34_tm_y+_q___pip_5160_1_53___block_40_dt_y;

// __block_1021
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1019
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1022
if (_t___block_1012_z_sel) begin
// __block_1023
// __block_1025
_d___pip_5160_1_53___stage___block_26_v_z = _q___pip_5160_1_53___stage___block_26_v_z+_q___pip_5160_1_53___stage___block_26_s_z;

_d___pip_5160_1_53___block_34_tm_z = _q___pip_5160_1_53___block_34_tm_z+_q___pip_5160_1_53___block_40_dt_z;

// __block_1026
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1024
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1027
// end of pipeline stage
_d__full_fsm___pip_5160_1_53 = 1;
_d__idx_fsm___pip_5160_1_53 = _t__stall_fsm___pip_5160_1_53 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_53 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 54
(* full_case *)
case (_q__idx_fsm___pip_5160_1_54)
1: begin
// __stage___block_1028
_t___stage___block_1028_tex = (_q___pip_5160_1_54___stage___block_26_v_x)^(_q___pip_5160_1_54___stage___block_26_v_y)^(_q___pip_5160_1_54___stage___block_26_v_z);

_t___stage___block_1028_vnum0 = {_q___pip_5160_1_54___stage___block_26_v_z[0+:2],_q___pip_5160_1_54___stage___block_26_v_y[0+:2],_q___pip_5160_1_54___stage___block_26_v_x[0+:2]};

_t___stage___block_1028_vnum1 = {_q___pip_5160_1_54___stage___block_26_v_z[2+:2],_q___pip_5160_1_54___stage___block_26_v_y[2+:2],_q___pip_5160_1_54___stage___block_26_v_x[2+:2]};

_t___stage___block_1028_vnum2 = {_q___pip_5160_1_54___stage___block_26_v_z[4+:2],_q___pip_5160_1_54___stage___block_26_v_y[4+:2],_q___pip_5160_1_54___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_54___stage___block_6_inside&_w_tile[_t___stage___block_1028_vnum0+:1]&_w_tile[_t___stage___block_1028_vnum1+:1]&_w_tile[_t___stage___block_1028_vnum2+:1]) begin
// __block_1029
// __block_1031
_d___pip_5160_1_54___stage___block_6_clr = _t___stage___block_1028_tex;

_d___pip_5160_1_54___stage___block_6_dist = 87;

_d___pip_5160_1_54___stage___block_6_inside = 1;

// __block_1032
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1030
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1033
_t___block_1033_cmp_yx = _q___pip_5160_1_54___block_34_tm_y-_q___pip_5160_1_54___block_34_tm_x;

_t___block_1033_cmp_zx = _q___pip_5160_1_54___block_34_tm_z-_q___pip_5160_1_54___block_34_tm_x;

_t___block_1033_cmp_zy = _q___pip_5160_1_54___block_34_tm_z-_q___pip_5160_1_54___block_34_tm_y;

_t___block_1033_x_sel = ~_t___block_1033_cmp_yx[20+:1]&&~_t___block_1033_cmp_zx[20+:1];

_t___block_1033_y_sel = _t___block_1033_cmp_yx[20+:1]&&~_t___block_1033_cmp_zy[20+:1];

_t___block_1033_z_sel = _t___block_1033_cmp_zx[20+:1]&&_t___block_1033_cmp_zy[20+:1];

if (_t___block_1033_x_sel) begin
// __block_1034
// __block_1036
_d___pip_5160_1_54___stage___block_26_v_x = _q___pip_5160_1_54___stage___block_26_v_x+_q___pip_5160_1_54___stage___block_26_s_x;

_d___pip_5160_1_54___block_34_tm_x = _q___pip_5160_1_54___block_34_tm_x+_q___pip_5160_1_54___block_40_dt_x;

// __block_1037
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1035
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1038
if (_t___block_1033_y_sel) begin
// __block_1039
// __block_1041
_d___pip_5160_1_54___stage___block_26_v_y = _q___pip_5160_1_54___stage___block_26_v_y+_q___pip_5160_1_54___stage___block_26_s_y;

_d___pip_5160_1_54___block_34_tm_y = _q___pip_5160_1_54___block_34_tm_y+_q___pip_5160_1_54___block_40_dt_y;

// __block_1042
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1040
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1043
if (_t___block_1033_z_sel) begin
// __block_1044
// __block_1046
_d___pip_5160_1_54___stage___block_26_v_z = _q___pip_5160_1_54___stage___block_26_v_z+_q___pip_5160_1_54___stage___block_26_s_z;

_d___pip_5160_1_54___block_34_tm_z = _q___pip_5160_1_54___block_34_tm_z+_q___pip_5160_1_54___block_40_dt_z;

// __block_1047
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1045
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1048
// end of pipeline stage
_d__full_fsm___pip_5160_1_54 = 1;
_d__idx_fsm___pip_5160_1_54 = _t__stall_fsm___pip_5160_1_54 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_54 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 55
(* full_case *)
case (_q__idx_fsm___pip_5160_1_55)
1: begin
// __stage___block_1049
_t___stage___block_1049_tex = (_q___pip_5160_1_55___stage___block_26_v_x)^(_q___pip_5160_1_55___stage___block_26_v_y)^(_q___pip_5160_1_55___stage___block_26_v_z);

_t___stage___block_1049_vnum0 = {_q___pip_5160_1_55___stage___block_26_v_z[0+:2],_q___pip_5160_1_55___stage___block_26_v_y[0+:2],_q___pip_5160_1_55___stage___block_26_v_x[0+:2]};

_t___stage___block_1049_vnum1 = {_q___pip_5160_1_55___stage___block_26_v_z[2+:2],_q___pip_5160_1_55___stage___block_26_v_y[2+:2],_q___pip_5160_1_55___stage___block_26_v_x[2+:2]};

_t___stage___block_1049_vnum2 = {_q___pip_5160_1_55___stage___block_26_v_z[4+:2],_q___pip_5160_1_55___stage___block_26_v_y[4+:2],_q___pip_5160_1_55___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_55___stage___block_6_inside&_w_tile[_t___stage___block_1049_vnum0+:1]&_w_tile[_t___stage___block_1049_vnum1+:1]&_w_tile[_t___stage___block_1049_vnum2+:1]) begin
// __block_1050
// __block_1052
_d___pip_5160_1_55___stage___block_6_clr = _t___stage___block_1049_tex;

_d___pip_5160_1_55___stage___block_6_dist = 89;

_d___pip_5160_1_55___stage___block_6_inside = 1;

// __block_1053
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1051
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1054
_t___block_1054_cmp_yx = _q___pip_5160_1_55___block_34_tm_y-_q___pip_5160_1_55___block_34_tm_x;

_t___block_1054_cmp_zx = _q___pip_5160_1_55___block_34_tm_z-_q___pip_5160_1_55___block_34_tm_x;

_t___block_1054_cmp_zy = _q___pip_5160_1_55___block_34_tm_z-_q___pip_5160_1_55___block_34_tm_y;

_t___block_1054_x_sel = ~_t___block_1054_cmp_yx[20+:1]&&~_t___block_1054_cmp_zx[20+:1];

_t___block_1054_y_sel = _t___block_1054_cmp_yx[20+:1]&&~_t___block_1054_cmp_zy[20+:1];

_t___block_1054_z_sel = _t___block_1054_cmp_zx[20+:1]&&_t___block_1054_cmp_zy[20+:1];

if (_t___block_1054_x_sel) begin
// __block_1055
// __block_1057
_d___pip_5160_1_55___stage___block_26_v_x = _q___pip_5160_1_55___stage___block_26_v_x+_q___pip_5160_1_55___stage___block_26_s_x;

_d___pip_5160_1_55___block_34_tm_x = _q___pip_5160_1_55___block_34_tm_x+_q___pip_5160_1_55___block_40_dt_x;

// __block_1058
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1056
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1059
if (_t___block_1054_y_sel) begin
// __block_1060
// __block_1062
_d___pip_5160_1_55___stage___block_26_v_y = _q___pip_5160_1_55___stage___block_26_v_y+_q___pip_5160_1_55___stage___block_26_s_y;

_d___pip_5160_1_55___block_34_tm_y = _q___pip_5160_1_55___block_34_tm_y+_q___pip_5160_1_55___block_40_dt_y;

// __block_1063
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1061
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1064
if (_t___block_1054_z_sel) begin
// __block_1065
// __block_1067
_d___pip_5160_1_55___stage___block_26_v_z = _q___pip_5160_1_55___stage___block_26_v_z+_q___pip_5160_1_55___stage___block_26_s_z;

_d___pip_5160_1_55___block_34_tm_z = _q___pip_5160_1_55___block_34_tm_z+_q___pip_5160_1_55___block_40_dt_z;

// __block_1068
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1066
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1069
// end of pipeline stage
_d__full_fsm___pip_5160_1_55 = 1;
_d__idx_fsm___pip_5160_1_55 = _t__stall_fsm___pip_5160_1_55 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_55 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 56
(* full_case *)
case (_q__idx_fsm___pip_5160_1_56)
1: begin
// __stage___block_1070
_t___stage___block_1070_tex = (_q___pip_5160_1_56___stage___block_26_v_x)^(_q___pip_5160_1_56___stage___block_26_v_y)^(_q___pip_5160_1_56___stage___block_26_v_z);

_t___stage___block_1070_vnum0 = {_q___pip_5160_1_56___stage___block_26_v_z[0+:2],_q___pip_5160_1_56___stage___block_26_v_y[0+:2],_q___pip_5160_1_56___stage___block_26_v_x[0+:2]};

_t___stage___block_1070_vnum1 = {_q___pip_5160_1_56___stage___block_26_v_z[2+:2],_q___pip_5160_1_56___stage___block_26_v_y[2+:2],_q___pip_5160_1_56___stage___block_26_v_x[2+:2]};

_t___stage___block_1070_vnum2 = {_q___pip_5160_1_56___stage___block_26_v_z[4+:2],_q___pip_5160_1_56___stage___block_26_v_y[4+:2],_q___pip_5160_1_56___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_56___stage___block_6_inside&_w_tile[_t___stage___block_1070_vnum0+:1]&_w_tile[_t___stage___block_1070_vnum1+:1]&_w_tile[_t___stage___block_1070_vnum2+:1]) begin
// __block_1071
// __block_1073
_d___pip_5160_1_56___stage___block_6_clr = _t___stage___block_1070_tex;

_d___pip_5160_1_56___stage___block_6_dist = 91;

_d___pip_5160_1_56___stage___block_6_inside = 1;

// __block_1074
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1072
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1075
_t___block_1075_cmp_yx = _q___pip_5160_1_56___block_34_tm_y-_q___pip_5160_1_56___block_34_tm_x;

_t___block_1075_cmp_zx = _q___pip_5160_1_56___block_34_tm_z-_q___pip_5160_1_56___block_34_tm_x;

_t___block_1075_cmp_zy = _q___pip_5160_1_56___block_34_tm_z-_q___pip_5160_1_56___block_34_tm_y;

_t___block_1075_x_sel = ~_t___block_1075_cmp_yx[20+:1]&&~_t___block_1075_cmp_zx[20+:1];

_t___block_1075_y_sel = _t___block_1075_cmp_yx[20+:1]&&~_t___block_1075_cmp_zy[20+:1];

_t___block_1075_z_sel = _t___block_1075_cmp_zx[20+:1]&&_t___block_1075_cmp_zy[20+:1];

if (_t___block_1075_x_sel) begin
// __block_1076
// __block_1078
_d___pip_5160_1_56___stage___block_26_v_x = _q___pip_5160_1_56___stage___block_26_v_x+_q___pip_5160_1_56___stage___block_26_s_x;

_d___pip_5160_1_56___block_34_tm_x = _q___pip_5160_1_56___block_34_tm_x+_q___pip_5160_1_56___block_40_dt_x;

// __block_1079
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1077
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1080
if (_t___block_1075_y_sel) begin
// __block_1081
// __block_1083
_d___pip_5160_1_56___stage___block_26_v_y = _q___pip_5160_1_56___stage___block_26_v_y+_q___pip_5160_1_56___stage___block_26_s_y;

_d___pip_5160_1_56___block_34_tm_y = _q___pip_5160_1_56___block_34_tm_y+_q___pip_5160_1_56___block_40_dt_y;

// __block_1084
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1082
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1085
if (_t___block_1075_z_sel) begin
// __block_1086
// __block_1088
_d___pip_5160_1_56___stage___block_26_v_z = _q___pip_5160_1_56___stage___block_26_v_z+_q___pip_5160_1_56___stage___block_26_s_z;

_d___pip_5160_1_56___block_34_tm_z = _q___pip_5160_1_56___block_34_tm_z+_q___pip_5160_1_56___block_40_dt_z;

// __block_1089
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1087
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1090
// end of pipeline stage
_d__full_fsm___pip_5160_1_56 = 1;
_d__idx_fsm___pip_5160_1_56 = _t__stall_fsm___pip_5160_1_56 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_56 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 57
(* full_case *)
case (_q__idx_fsm___pip_5160_1_57)
1: begin
// __stage___block_1091
_t___stage___block_1091_tex = (_q___pip_5160_1_57___stage___block_26_v_x)^(_q___pip_5160_1_57___stage___block_26_v_y)^(_q___pip_5160_1_57___stage___block_26_v_z);

_t___stage___block_1091_vnum0 = {_q___pip_5160_1_57___stage___block_26_v_z[0+:2],_q___pip_5160_1_57___stage___block_26_v_y[0+:2],_q___pip_5160_1_57___stage___block_26_v_x[0+:2]};

_t___stage___block_1091_vnum1 = {_q___pip_5160_1_57___stage___block_26_v_z[2+:2],_q___pip_5160_1_57___stage___block_26_v_y[2+:2],_q___pip_5160_1_57___stage___block_26_v_x[2+:2]};

_t___stage___block_1091_vnum2 = {_q___pip_5160_1_57___stage___block_26_v_z[4+:2],_q___pip_5160_1_57___stage___block_26_v_y[4+:2],_q___pip_5160_1_57___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_57___stage___block_6_inside&_w_tile[_t___stage___block_1091_vnum0+:1]&_w_tile[_t___stage___block_1091_vnum1+:1]&_w_tile[_t___stage___block_1091_vnum2+:1]) begin
// __block_1092
// __block_1094
_d___pip_5160_1_57___stage___block_6_clr = _t___stage___block_1091_tex;

_d___pip_5160_1_57___stage___block_6_dist = 93;

_d___pip_5160_1_57___stage___block_6_inside = 1;

// __block_1095
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1093
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1096
_t___block_1096_cmp_yx = _q___pip_5160_1_57___block_34_tm_y-_q___pip_5160_1_57___block_34_tm_x;

_t___block_1096_cmp_zx = _q___pip_5160_1_57___block_34_tm_z-_q___pip_5160_1_57___block_34_tm_x;

_t___block_1096_cmp_zy = _q___pip_5160_1_57___block_34_tm_z-_q___pip_5160_1_57___block_34_tm_y;

_t___block_1096_x_sel = ~_t___block_1096_cmp_yx[20+:1]&&~_t___block_1096_cmp_zx[20+:1];

_t___block_1096_y_sel = _t___block_1096_cmp_yx[20+:1]&&~_t___block_1096_cmp_zy[20+:1];

_t___block_1096_z_sel = _t___block_1096_cmp_zx[20+:1]&&_t___block_1096_cmp_zy[20+:1];

if (_t___block_1096_x_sel) begin
// __block_1097
// __block_1099
_d___pip_5160_1_57___stage___block_26_v_x = _q___pip_5160_1_57___stage___block_26_v_x+_q___pip_5160_1_57___stage___block_26_s_x;

_d___pip_5160_1_57___block_34_tm_x = _q___pip_5160_1_57___block_34_tm_x+_q___pip_5160_1_57___block_40_dt_x;

// __block_1100
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1098
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1101
if (_t___block_1096_y_sel) begin
// __block_1102
// __block_1104
_d___pip_5160_1_57___stage___block_26_v_y = _q___pip_5160_1_57___stage___block_26_v_y+_q___pip_5160_1_57___stage___block_26_s_y;

_d___pip_5160_1_57___block_34_tm_y = _q___pip_5160_1_57___block_34_tm_y+_q___pip_5160_1_57___block_40_dt_y;

// __block_1105
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1103
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1106
if (_t___block_1096_z_sel) begin
// __block_1107
// __block_1109
_d___pip_5160_1_57___stage___block_26_v_z = _q___pip_5160_1_57___stage___block_26_v_z+_q___pip_5160_1_57___stage___block_26_s_z;

_d___pip_5160_1_57___block_34_tm_z = _q___pip_5160_1_57___block_34_tm_z+_q___pip_5160_1_57___block_40_dt_z;

// __block_1110
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1108
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1111
// end of pipeline stage
_d__full_fsm___pip_5160_1_57 = 1;
_d__idx_fsm___pip_5160_1_57 = _t__stall_fsm___pip_5160_1_57 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_57 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 58
(* full_case *)
case (_q__idx_fsm___pip_5160_1_58)
1: begin
// __stage___block_1112
_t___stage___block_1112_tex = (_q___pip_5160_1_58___stage___block_26_v_x)^(_q___pip_5160_1_58___stage___block_26_v_y)^(_q___pip_5160_1_58___stage___block_26_v_z);

_t___stage___block_1112_vnum0 = {_q___pip_5160_1_58___stage___block_26_v_z[0+:2],_q___pip_5160_1_58___stage___block_26_v_y[0+:2],_q___pip_5160_1_58___stage___block_26_v_x[0+:2]};

_t___stage___block_1112_vnum1 = {_q___pip_5160_1_58___stage___block_26_v_z[2+:2],_q___pip_5160_1_58___stage___block_26_v_y[2+:2],_q___pip_5160_1_58___stage___block_26_v_x[2+:2]};

_t___stage___block_1112_vnum2 = {_q___pip_5160_1_58___stage___block_26_v_z[4+:2],_q___pip_5160_1_58___stage___block_26_v_y[4+:2],_q___pip_5160_1_58___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_58___stage___block_6_inside&_w_tile[_t___stage___block_1112_vnum0+:1]&_w_tile[_t___stage___block_1112_vnum1+:1]&_w_tile[_t___stage___block_1112_vnum2+:1]) begin
// __block_1113
// __block_1115
_d___pip_5160_1_58___stage___block_6_clr = _t___stage___block_1112_tex;

_d___pip_5160_1_58___stage___block_6_dist = 95;

_d___pip_5160_1_58___stage___block_6_inside = 1;

// __block_1116
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1114
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1117
_t___block_1117_cmp_yx = _q___pip_5160_1_58___block_34_tm_y-_q___pip_5160_1_58___block_34_tm_x;

_t___block_1117_cmp_zx = _q___pip_5160_1_58___block_34_tm_z-_q___pip_5160_1_58___block_34_tm_x;

_t___block_1117_cmp_zy = _q___pip_5160_1_58___block_34_tm_z-_q___pip_5160_1_58___block_34_tm_y;

_t___block_1117_x_sel = ~_t___block_1117_cmp_yx[20+:1]&&~_t___block_1117_cmp_zx[20+:1];

_t___block_1117_y_sel = _t___block_1117_cmp_yx[20+:1]&&~_t___block_1117_cmp_zy[20+:1];

_t___block_1117_z_sel = _t___block_1117_cmp_zx[20+:1]&&_t___block_1117_cmp_zy[20+:1];

if (_t___block_1117_x_sel) begin
// __block_1118
// __block_1120
_d___pip_5160_1_58___stage___block_26_v_x = _q___pip_5160_1_58___stage___block_26_v_x+_q___pip_5160_1_58___stage___block_26_s_x;

_d___pip_5160_1_58___block_34_tm_x = _q___pip_5160_1_58___block_34_tm_x+_q___pip_5160_1_58___block_40_dt_x;

// __block_1121
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1119
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1122
if (_t___block_1117_y_sel) begin
// __block_1123
// __block_1125
_d___pip_5160_1_58___stage___block_26_v_y = _q___pip_5160_1_58___stage___block_26_v_y+_q___pip_5160_1_58___stage___block_26_s_y;

_d___pip_5160_1_58___block_34_tm_y = _q___pip_5160_1_58___block_34_tm_y+_q___pip_5160_1_58___block_40_dt_y;

// __block_1126
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1124
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1127
if (_t___block_1117_z_sel) begin
// __block_1128
// __block_1130
_d___pip_5160_1_58___stage___block_26_v_z = _q___pip_5160_1_58___stage___block_26_v_z+_q___pip_5160_1_58___stage___block_26_s_z;

_d___pip_5160_1_58___block_34_tm_z = _q___pip_5160_1_58___block_34_tm_z+_q___pip_5160_1_58___block_40_dt_z;

// __block_1131
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1129
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1132
// end of pipeline stage
_d__full_fsm___pip_5160_1_58 = 1;
_d__idx_fsm___pip_5160_1_58 = _t__stall_fsm___pip_5160_1_58 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_58 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 59
(* full_case *)
case (_q__idx_fsm___pip_5160_1_59)
1: begin
// __stage___block_1133
_t___stage___block_1133_tex = (_q___pip_5160_1_59___stage___block_26_v_x)^(_q___pip_5160_1_59___stage___block_26_v_y)^(_q___pip_5160_1_59___stage___block_26_v_z);

_t___stage___block_1133_vnum0 = {_q___pip_5160_1_59___stage___block_26_v_z[0+:2],_q___pip_5160_1_59___stage___block_26_v_y[0+:2],_q___pip_5160_1_59___stage___block_26_v_x[0+:2]};

_t___stage___block_1133_vnum1 = {_q___pip_5160_1_59___stage___block_26_v_z[2+:2],_q___pip_5160_1_59___stage___block_26_v_y[2+:2],_q___pip_5160_1_59___stage___block_26_v_x[2+:2]};

_t___stage___block_1133_vnum2 = {_q___pip_5160_1_59___stage___block_26_v_z[4+:2],_q___pip_5160_1_59___stage___block_26_v_y[4+:2],_q___pip_5160_1_59___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_59___stage___block_6_inside&_w_tile[_t___stage___block_1133_vnum0+:1]&_w_tile[_t___stage___block_1133_vnum1+:1]&_w_tile[_t___stage___block_1133_vnum2+:1]) begin
// __block_1134
// __block_1136
_d___pip_5160_1_59___stage___block_6_clr = _t___stage___block_1133_tex;

_d___pip_5160_1_59___stage___block_6_dist = 97;

_d___pip_5160_1_59___stage___block_6_inside = 1;

// __block_1137
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1135
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1138
_t___block_1138_cmp_yx = _q___pip_5160_1_59___block_34_tm_y-_q___pip_5160_1_59___block_34_tm_x;

_t___block_1138_cmp_zx = _q___pip_5160_1_59___block_34_tm_z-_q___pip_5160_1_59___block_34_tm_x;

_t___block_1138_cmp_zy = _q___pip_5160_1_59___block_34_tm_z-_q___pip_5160_1_59___block_34_tm_y;

_t___block_1138_x_sel = ~_t___block_1138_cmp_yx[20+:1]&&~_t___block_1138_cmp_zx[20+:1];

_t___block_1138_y_sel = _t___block_1138_cmp_yx[20+:1]&&~_t___block_1138_cmp_zy[20+:1];

_t___block_1138_z_sel = _t___block_1138_cmp_zx[20+:1]&&_t___block_1138_cmp_zy[20+:1];

if (_t___block_1138_x_sel) begin
// __block_1139
// __block_1141
_d___pip_5160_1_59___stage___block_26_v_x = _q___pip_5160_1_59___stage___block_26_v_x+_q___pip_5160_1_59___stage___block_26_s_x;

_d___pip_5160_1_59___block_34_tm_x = _q___pip_5160_1_59___block_34_tm_x+_q___pip_5160_1_59___block_40_dt_x;

// __block_1142
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1140
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1143
if (_t___block_1138_y_sel) begin
// __block_1144
// __block_1146
_d___pip_5160_1_59___stage___block_26_v_y = _q___pip_5160_1_59___stage___block_26_v_y+_q___pip_5160_1_59___stage___block_26_s_y;

_d___pip_5160_1_59___block_34_tm_y = _q___pip_5160_1_59___block_34_tm_y+_q___pip_5160_1_59___block_40_dt_y;

// __block_1147
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1145
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1148
if (_t___block_1138_z_sel) begin
// __block_1149
// __block_1151
_d___pip_5160_1_59___stage___block_26_v_z = _q___pip_5160_1_59___stage___block_26_v_z+_q___pip_5160_1_59___stage___block_26_s_z;

_d___pip_5160_1_59___block_34_tm_z = _q___pip_5160_1_59___block_34_tm_z+_q___pip_5160_1_59___block_40_dt_z;

// __block_1152
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1150
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1153
// end of pipeline stage
_d__full_fsm___pip_5160_1_59 = 1;
_d__idx_fsm___pip_5160_1_59 = _t__stall_fsm___pip_5160_1_59 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_59 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 60
(* full_case *)
case (_q__idx_fsm___pip_5160_1_60)
1: begin
// __stage___block_1154
_t___stage___block_1154_tex = (_q___pip_5160_1_60___stage___block_26_v_x)^(_q___pip_5160_1_60___stage___block_26_v_y)^(_q___pip_5160_1_60___stage___block_26_v_z);

_t___stage___block_1154_vnum0 = {_q___pip_5160_1_60___stage___block_26_v_z[0+:2],_q___pip_5160_1_60___stage___block_26_v_y[0+:2],_q___pip_5160_1_60___stage___block_26_v_x[0+:2]};

_t___stage___block_1154_vnum1 = {_q___pip_5160_1_60___stage___block_26_v_z[2+:2],_q___pip_5160_1_60___stage___block_26_v_y[2+:2],_q___pip_5160_1_60___stage___block_26_v_x[2+:2]};

_t___stage___block_1154_vnum2 = {_q___pip_5160_1_60___stage___block_26_v_z[4+:2],_q___pip_5160_1_60___stage___block_26_v_y[4+:2],_q___pip_5160_1_60___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_60___stage___block_6_inside&_w_tile[_t___stage___block_1154_vnum0+:1]&_w_tile[_t___stage___block_1154_vnum1+:1]&_w_tile[_t___stage___block_1154_vnum2+:1]) begin
// __block_1155
// __block_1157
_d___pip_5160_1_60___stage___block_6_clr = _t___stage___block_1154_tex;

_d___pip_5160_1_60___stage___block_6_dist = 98;

_d___pip_5160_1_60___stage___block_6_inside = 1;

// __block_1158
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1156
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1159
_t___block_1159_cmp_yx = _q___pip_5160_1_60___block_34_tm_y-_q___pip_5160_1_60___block_34_tm_x;

_t___block_1159_cmp_zx = _q___pip_5160_1_60___block_34_tm_z-_q___pip_5160_1_60___block_34_tm_x;

_t___block_1159_cmp_zy = _q___pip_5160_1_60___block_34_tm_z-_q___pip_5160_1_60___block_34_tm_y;

_t___block_1159_x_sel = ~_t___block_1159_cmp_yx[20+:1]&&~_t___block_1159_cmp_zx[20+:1];

_t___block_1159_y_sel = _t___block_1159_cmp_yx[20+:1]&&~_t___block_1159_cmp_zy[20+:1];

_t___block_1159_z_sel = _t___block_1159_cmp_zx[20+:1]&&_t___block_1159_cmp_zy[20+:1];

if (_t___block_1159_x_sel) begin
// __block_1160
// __block_1162
_d___pip_5160_1_60___stage___block_26_v_x = _q___pip_5160_1_60___stage___block_26_v_x+_q___pip_5160_1_60___stage___block_26_s_x;

_d___pip_5160_1_60___block_34_tm_x = _q___pip_5160_1_60___block_34_tm_x+_q___pip_5160_1_60___block_40_dt_x;

// __block_1163
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1161
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1164
if (_t___block_1159_y_sel) begin
// __block_1165
// __block_1167
_d___pip_5160_1_60___stage___block_26_v_y = _q___pip_5160_1_60___stage___block_26_v_y+_q___pip_5160_1_60___stage___block_26_s_y;

_d___pip_5160_1_60___block_34_tm_y = _q___pip_5160_1_60___block_34_tm_y+_q___pip_5160_1_60___block_40_dt_y;

// __block_1168
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1166
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1169
if (_t___block_1159_z_sel) begin
// __block_1170
// __block_1172
_d___pip_5160_1_60___stage___block_26_v_z = _q___pip_5160_1_60___stage___block_26_v_z+_q___pip_5160_1_60___stage___block_26_s_z;

_d___pip_5160_1_60___block_34_tm_z = _q___pip_5160_1_60___block_34_tm_z+_q___pip_5160_1_60___block_40_dt_z;

// __block_1173
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1171
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1174
// end of pipeline stage
_d__full_fsm___pip_5160_1_60 = 1;
_d__idx_fsm___pip_5160_1_60 = _t__stall_fsm___pip_5160_1_60 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_60 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 61
(* full_case *)
case (_q__idx_fsm___pip_5160_1_61)
1: begin
// __stage___block_1175
_t___stage___block_1175_tex = (_q___pip_5160_1_61___stage___block_26_v_x)^(_q___pip_5160_1_61___stage___block_26_v_y)^(_q___pip_5160_1_61___stage___block_26_v_z);

_t___stage___block_1175_vnum0 = {_q___pip_5160_1_61___stage___block_26_v_z[0+:2],_q___pip_5160_1_61___stage___block_26_v_y[0+:2],_q___pip_5160_1_61___stage___block_26_v_x[0+:2]};

_t___stage___block_1175_vnum1 = {_q___pip_5160_1_61___stage___block_26_v_z[2+:2],_q___pip_5160_1_61___stage___block_26_v_y[2+:2],_q___pip_5160_1_61___stage___block_26_v_x[2+:2]};

_t___stage___block_1175_vnum2 = {_q___pip_5160_1_61___stage___block_26_v_z[4+:2],_q___pip_5160_1_61___stage___block_26_v_y[4+:2],_q___pip_5160_1_61___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_61___stage___block_6_inside&_w_tile[_t___stage___block_1175_vnum0+:1]&_w_tile[_t___stage___block_1175_vnum1+:1]&_w_tile[_t___stage___block_1175_vnum2+:1]) begin
// __block_1176
// __block_1178
_d___pip_5160_1_61___stage___block_6_clr = _t___stage___block_1175_tex;

_d___pip_5160_1_61___stage___block_6_dist = 100;

_d___pip_5160_1_61___stage___block_6_inside = 1;

// __block_1179
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1177
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1180
_t___block_1180_cmp_yx = _q___pip_5160_1_61___block_34_tm_y-_q___pip_5160_1_61___block_34_tm_x;

_t___block_1180_cmp_zx = _q___pip_5160_1_61___block_34_tm_z-_q___pip_5160_1_61___block_34_tm_x;

_t___block_1180_cmp_zy = _q___pip_5160_1_61___block_34_tm_z-_q___pip_5160_1_61___block_34_tm_y;

_t___block_1180_x_sel = ~_t___block_1180_cmp_yx[20+:1]&&~_t___block_1180_cmp_zx[20+:1];

_t___block_1180_y_sel = _t___block_1180_cmp_yx[20+:1]&&~_t___block_1180_cmp_zy[20+:1];

_t___block_1180_z_sel = _t___block_1180_cmp_zx[20+:1]&&_t___block_1180_cmp_zy[20+:1];

if (_t___block_1180_x_sel) begin
// __block_1181
// __block_1183
_d___pip_5160_1_61___stage___block_26_v_x = _q___pip_5160_1_61___stage___block_26_v_x+_q___pip_5160_1_61___stage___block_26_s_x;

_d___pip_5160_1_61___block_34_tm_x = _q___pip_5160_1_61___block_34_tm_x+_q___pip_5160_1_61___block_40_dt_x;

// __block_1184
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1182
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1185
if (_t___block_1180_y_sel) begin
// __block_1186
// __block_1188
_d___pip_5160_1_61___stage___block_26_v_y = _q___pip_5160_1_61___stage___block_26_v_y+_q___pip_5160_1_61___stage___block_26_s_y;

_d___pip_5160_1_61___block_34_tm_y = _q___pip_5160_1_61___block_34_tm_y+_q___pip_5160_1_61___block_40_dt_y;

// __block_1189
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1187
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1190
if (_t___block_1180_z_sel) begin
// __block_1191
// __block_1193
_d___pip_5160_1_61___stage___block_26_v_z = _q___pip_5160_1_61___stage___block_26_v_z+_q___pip_5160_1_61___stage___block_26_s_z;

_d___pip_5160_1_61___block_34_tm_z = _q___pip_5160_1_61___block_34_tm_z+_q___pip_5160_1_61___block_40_dt_z;

// __block_1194
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1192
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1195
// end of pipeline stage
_d__full_fsm___pip_5160_1_61 = 1;
_d__idx_fsm___pip_5160_1_61 = _t__stall_fsm___pip_5160_1_61 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_61 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 62
(* full_case *)
case (_q__idx_fsm___pip_5160_1_62)
1: begin
// __stage___block_1196
_t___stage___block_1196_tex = (_q___pip_5160_1_62___stage___block_26_v_x)^(_q___pip_5160_1_62___stage___block_26_v_y)^(_q___pip_5160_1_62___stage___block_26_v_z);

_t___stage___block_1196_vnum0 = {_q___pip_5160_1_62___stage___block_26_v_z[0+:2],_q___pip_5160_1_62___stage___block_26_v_y[0+:2],_q___pip_5160_1_62___stage___block_26_v_x[0+:2]};

_t___stage___block_1196_vnum1 = {_q___pip_5160_1_62___stage___block_26_v_z[2+:2],_q___pip_5160_1_62___stage___block_26_v_y[2+:2],_q___pip_5160_1_62___stage___block_26_v_x[2+:2]};

_t___stage___block_1196_vnum2 = {_q___pip_5160_1_62___stage___block_26_v_z[4+:2],_q___pip_5160_1_62___stage___block_26_v_y[4+:2],_q___pip_5160_1_62___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_62___stage___block_6_inside&_w_tile[_t___stage___block_1196_vnum0+:1]&_w_tile[_t___stage___block_1196_vnum1+:1]&_w_tile[_t___stage___block_1196_vnum2+:1]) begin
// __block_1197
// __block_1199
_d___pip_5160_1_62___stage___block_6_clr = _t___stage___block_1196_tex;

_d___pip_5160_1_62___stage___block_6_dist = 102;

_d___pip_5160_1_62___stage___block_6_inside = 1;

// __block_1200
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1198
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1201
_t___block_1201_cmp_yx = _q___pip_5160_1_62___block_34_tm_y-_q___pip_5160_1_62___block_34_tm_x;

_t___block_1201_cmp_zx = _q___pip_5160_1_62___block_34_tm_z-_q___pip_5160_1_62___block_34_tm_x;

_t___block_1201_cmp_zy = _q___pip_5160_1_62___block_34_tm_z-_q___pip_5160_1_62___block_34_tm_y;

_t___block_1201_x_sel = ~_t___block_1201_cmp_yx[20+:1]&&~_t___block_1201_cmp_zx[20+:1];

_t___block_1201_y_sel = _t___block_1201_cmp_yx[20+:1]&&~_t___block_1201_cmp_zy[20+:1];

_t___block_1201_z_sel = _t___block_1201_cmp_zx[20+:1]&&_t___block_1201_cmp_zy[20+:1];

if (_t___block_1201_x_sel) begin
// __block_1202
// __block_1204
_d___pip_5160_1_62___stage___block_26_v_x = _q___pip_5160_1_62___stage___block_26_v_x+_q___pip_5160_1_62___stage___block_26_s_x;

_d___pip_5160_1_62___block_34_tm_x = _q___pip_5160_1_62___block_34_tm_x+_q___pip_5160_1_62___block_40_dt_x;

// __block_1205
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1203
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1206
if (_t___block_1201_y_sel) begin
// __block_1207
// __block_1209
_d___pip_5160_1_62___stage___block_26_v_y = _q___pip_5160_1_62___stage___block_26_v_y+_q___pip_5160_1_62___stage___block_26_s_y;

_d___pip_5160_1_62___block_34_tm_y = _q___pip_5160_1_62___block_34_tm_y+_q___pip_5160_1_62___block_40_dt_y;

// __block_1210
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1208
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1211
if (_t___block_1201_z_sel) begin
// __block_1212
// __block_1214
_d___pip_5160_1_62___stage___block_26_v_z = _q___pip_5160_1_62___stage___block_26_v_z+_q___pip_5160_1_62___stage___block_26_s_z;

_d___pip_5160_1_62___block_34_tm_z = _q___pip_5160_1_62___block_34_tm_z+_q___pip_5160_1_62___block_40_dt_z;

// __block_1215
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1213
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1216
// end of pipeline stage
_d__full_fsm___pip_5160_1_62 = 1;
_d__idx_fsm___pip_5160_1_62 = _t__stall_fsm___pip_5160_1_62 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_62 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 63
(* full_case *)
case (_q__idx_fsm___pip_5160_1_63)
1: begin
// __stage___block_1217
_t___stage___block_1217_tex = (_q___pip_5160_1_63___stage___block_26_v_x)^(_q___pip_5160_1_63___stage___block_26_v_y)^(_q___pip_5160_1_63___stage___block_26_v_z);

_t___stage___block_1217_vnum0 = {_q___pip_5160_1_63___stage___block_26_v_z[0+:2],_q___pip_5160_1_63___stage___block_26_v_y[0+:2],_q___pip_5160_1_63___stage___block_26_v_x[0+:2]};

_t___stage___block_1217_vnum1 = {_q___pip_5160_1_63___stage___block_26_v_z[2+:2],_q___pip_5160_1_63___stage___block_26_v_y[2+:2],_q___pip_5160_1_63___stage___block_26_v_x[2+:2]};

_t___stage___block_1217_vnum2 = {_q___pip_5160_1_63___stage___block_26_v_z[4+:2],_q___pip_5160_1_63___stage___block_26_v_y[4+:2],_q___pip_5160_1_63___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_63___stage___block_6_inside&_w_tile[_t___stage___block_1217_vnum0+:1]&_w_tile[_t___stage___block_1217_vnum1+:1]&_w_tile[_t___stage___block_1217_vnum2+:1]) begin
// __block_1218
// __block_1220
_d___pip_5160_1_63___stage___block_6_clr = _t___stage___block_1217_tex;

_d___pip_5160_1_63___stage___block_6_dist = 104;

_d___pip_5160_1_63___stage___block_6_inside = 1;

// __block_1221
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1219
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1222
_t___block_1222_cmp_yx = _q___pip_5160_1_63___block_34_tm_y-_q___pip_5160_1_63___block_34_tm_x;

_t___block_1222_cmp_zx = _q___pip_5160_1_63___block_34_tm_z-_q___pip_5160_1_63___block_34_tm_x;

_t___block_1222_cmp_zy = _q___pip_5160_1_63___block_34_tm_z-_q___pip_5160_1_63___block_34_tm_y;

_t___block_1222_x_sel = ~_t___block_1222_cmp_yx[20+:1]&&~_t___block_1222_cmp_zx[20+:1];

_t___block_1222_y_sel = _t___block_1222_cmp_yx[20+:1]&&~_t___block_1222_cmp_zy[20+:1];

_t___block_1222_z_sel = _t___block_1222_cmp_zx[20+:1]&&_t___block_1222_cmp_zy[20+:1];

if (_t___block_1222_x_sel) begin
// __block_1223
// __block_1225
_d___pip_5160_1_63___stage___block_26_v_x = _q___pip_5160_1_63___stage___block_26_v_x+_q___pip_5160_1_63___stage___block_26_s_x;

_d___pip_5160_1_63___block_34_tm_x = _q___pip_5160_1_63___block_34_tm_x+_q___pip_5160_1_63___block_40_dt_x;

// __block_1226
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1224
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1227
if (_t___block_1222_y_sel) begin
// __block_1228
// __block_1230
_d___pip_5160_1_63___stage___block_26_v_y = _q___pip_5160_1_63___stage___block_26_v_y+_q___pip_5160_1_63___stage___block_26_s_y;

_d___pip_5160_1_63___block_34_tm_y = _q___pip_5160_1_63___block_34_tm_y+_q___pip_5160_1_63___block_40_dt_y;

// __block_1231
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1229
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1232
if (_t___block_1222_z_sel) begin
// __block_1233
// __block_1235
_d___pip_5160_1_63___stage___block_26_v_z = _q___pip_5160_1_63___stage___block_26_v_z+_q___pip_5160_1_63___stage___block_26_s_z;

_d___pip_5160_1_63___block_34_tm_z = _q___pip_5160_1_63___block_34_tm_z+_q___pip_5160_1_63___block_40_dt_z;

// __block_1236
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1234
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1237
// end of pipeline stage
_d__full_fsm___pip_5160_1_63 = 1;
_d__idx_fsm___pip_5160_1_63 = _t__stall_fsm___pip_5160_1_63 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_63 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 64
(* full_case *)
case (_q__idx_fsm___pip_5160_1_64)
1: begin
// __stage___block_1238
_t___stage___block_1238_tex = (_q___pip_5160_1_64___stage___block_26_v_x)^(_q___pip_5160_1_64___stage___block_26_v_y)^(_q___pip_5160_1_64___stage___block_26_v_z);

_t___stage___block_1238_vnum0 = {_q___pip_5160_1_64___stage___block_26_v_z[0+:2],_q___pip_5160_1_64___stage___block_26_v_y[0+:2],_q___pip_5160_1_64___stage___block_26_v_x[0+:2]};

_t___stage___block_1238_vnum1 = {_q___pip_5160_1_64___stage___block_26_v_z[2+:2],_q___pip_5160_1_64___stage___block_26_v_y[2+:2],_q___pip_5160_1_64___stage___block_26_v_x[2+:2]};

_t___stage___block_1238_vnum2 = {_q___pip_5160_1_64___stage___block_26_v_z[4+:2],_q___pip_5160_1_64___stage___block_26_v_y[4+:2],_q___pip_5160_1_64___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_64___stage___block_6_inside&_w_tile[_t___stage___block_1238_vnum0+:1]&_w_tile[_t___stage___block_1238_vnum1+:1]&_w_tile[_t___stage___block_1238_vnum2+:1]) begin
// __block_1239
// __block_1241
_d___pip_5160_1_64___stage___block_6_clr = _t___stage___block_1238_tex;

_d___pip_5160_1_64___stage___block_6_dist = 106;

_d___pip_5160_1_64___stage___block_6_inside = 1;

// __block_1242
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1240
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1243
_t___block_1243_cmp_yx = _q___pip_5160_1_64___block_34_tm_y-_q___pip_5160_1_64___block_34_tm_x;

_t___block_1243_cmp_zx = _q___pip_5160_1_64___block_34_tm_z-_q___pip_5160_1_64___block_34_tm_x;

_t___block_1243_cmp_zy = _q___pip_5160_1_64___block_34_tm_z-_q___pip_5160_1_64___block_34_tm_y;

_t___block_1243_x_sel = ~_t___block_1243_cmp_yx[20+:1]&&~_t___block_1243_cmp_zx[20+:1];

_t___block_1243_y_sel = _t___block_1243_cmp_yx[20+:1]&&~_t___block_1243_cmp_zy[20+:1];

_t___block_1243_z_sel = _t___block_1243_cmp_zx[20+:1]&&_t___block_1243_cmp_zy[20+:1];

if (_t___block_1243_x_sel) begin
// __block_1244
// __block_1246
_d___pip_5160_1_64___stage___block_26_v_x = _q___pip_5160_1_64___stage___block_26_v_x+_q___pip_5160_1_64___stage___block_26_s_x;

_d___pip_5160_1_64___block_34_tm_x = _q___pip_5160_1_64___block_34_tm_x+_q___pip_5160_1_64___block_40_dt_x;

// __block_1247
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1245
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1248
if (_t___block_1243_y_sel) begin
// __block_1249
// __block_1251
_d___pip_5160_1_64___stage___block_26_v_y = _q___pip_5160_1_64___stage___block_26_v_y+_q___pip_5160_1_64___stage___block_26_s_y;

_d___pip_5160_1_64___block_34_tm_y = _q___pip_5160_1_64___block_34_tm_y+_q___pip_5160_1_64___block_40_dt_y;

// __block_1252
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1250
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1253
if (_t___block_1243_z_sel) begin
// __block_1254
// __block_1256
_d___pip_5160_1_64___stage___block_26_v_z = _q___pip_5160_1_64___stage___block_26_v_z+_q___pip_5160_1_64___stage___block_26_s_z;

_d___pip_5160_1_64___block_34_tm_z = _q___pip_5160_1_64___block_34_tm_z+_q___pip_5160_1_64___block_40_dt_z;

// __block_1257
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1255
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1258
// end of pipeline stage
_d__full_fsm___pip_5160_1_64 = 1;
_d__idx_fsm___pip_5160_1_64 = _t__stall_fsm___pip_5160_1_64 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_64 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 65
(* full_case *)
case (_q__idx_fsm___pip_5160_1_65)
1: begin
// __stage___block_1259
_t___stage___block_1259_tex = (_q___pip_5160_1_65___stage___block_26_v_x)^(_q___pip_5160_1_65___stage___block_26_v_y)^(_q___pip_5160_1_65___stage___block_26_v_z);

_t___stage___block_1259_vnum0 = {_q___pip_5160_1_65___stage___block_26_v_z[0+:2],_q___pip_5160_1_65___stage___block_26_v_y[0+:2],_q___pip_5160_1_65___stage___block_26_v_x[0+:2]};

_t___stage___block_1259_vnum1 = {_q___pip_5160_1_65___stage___block_26_v_z[2+:2],_q___pip_5160_1_65___stage___block_26_v_y[2+:2],_q___pip_5160_1_65___stage___block_26_v_x[2+:2]};

_t___stage___block_1259_vnum2 = {_q___pip_5160_1_65___stage___block_26_v_z[4+:2],_q___pip_5160_1_65___stage___block_26_v_y[4+:2],_q___pip_5160_1_65___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_65___stage___block_6_inside&_w_tile[_t___stage___block_1259_vnum0+:1]&_w_tile[_t___stage___block_1259_vnum1+:1]&_w_tile[_t___stage___block_1259_vnum2+:1]) begin
// __block_1260
// __block_1262
_d___pip_5160_1_65___stage___block_6_clr = _t___stage___block_1259_tex;

_d___pip_5160_1_65___stage___block_6_dist = 108;

_d___pip_5160_1_65___stage___block_6_inside = 1;

// __block_1263
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1261
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1264
_t___block_1264_cmp_yx = _q___pip_5160_1_65___block_34_tm_y-_q___pip_5160_1_65___block_34_tm_x;

_t___block_1264_cmp_zx = _q___pip_5160_1_65___block_34_tm_z-_q___pip_5160_1_65___block_34_tm_x;

_t___block_1264_cmp_zy = _q___pip_5160_1_65___block_34_tm_z-_q___pip_5160_1_65___block_34_tm_y;

_t___block_1264_x_sel = ~_t___block_1264_cmp_yx[20+:1]&&~_t___block_1264_cmp_zx[20+:1];

_t___block_1264_y_sel = _t___block_1264_cmp_yx[20+:1]&&~_t___block_1264_cmp_zy[20+:1];

_t___block_1264_z_sel = _t___block_1264_cmp_zx[20+:1]&&_t___block_1264_cmp_zy[20+:1];

if (_t___block_1264_x_sel) begin
// __block_1265
// __block_1267
_d___pip_5160_1_65___stage___block_26_v_x = _q___pip_5160_1_65___stage___block_26_v_x+_q___pip_5160_1_65___stage___block_26_s_x;

_d___pip_5160_1_65___block_34_tm_x = _q___pip_5160_1_65___block_34_tm_x+_q___pip_5160_1_65___block_40_dt_x;

// __block_1268
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1266
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1269
if (_t___block_1264_y_sel) begin
// __block_1270
// __block_1272
_d___pip_5160_1_65___stage___block_26_v_y = _q___pip_5160_1_65___stage___block_26_v_y+_q___pip_5160_1_65___stage___block_26_s_y;

_d___pip_5160_1_65___block_34_tm_y = _q___pip_5160_1_65___block_34_tm_y+_q___pip_5160_1_65___block_40_dt_y;

// __block_1273
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1271
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1274
if (_t___block_1264_z_sel) begin
// __block_1275
// __block_1277
_d___pip_5160_1_65___stage___block_26_v_z = _q___pip_5160_1_65___stage___block_26_v_z+_q___pip_5160_1_65___stage___block_26_s_z;

_d___pip_5160_1_65___block_34_tm_z = _q___pip_5160_1_65___block_34_tm_z+_q___pip_5160_1_65___block_40_dt_z;

// __block_1278
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1276
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1279
// end of pipeline stage
_d__full_fsm___pip_5160_1_65 = 1;
_d__idx_fsm___pip_5160_1_65 = _t__stall_fsm___pip_5160_1_65 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_65 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 66
(* full_case *)
case (_q__idx_fsm___pip_5160_1_66)
1: begin
// __stage___block_1280
_t___stage___block_1280_tex = (_q___pip_5160_1_66___stage___block_26_v_x)^(_q___pip_5160_1_66___stage___block_26_v_y)^(_q___pip_5160_1_66___stage___block_26_v_z);

_t___stage___block_1280_vnum0 = {_q___pip_5160_1_66___stage___block_26_v_z[0+:2],_q___pip_5160_1_66___stage___block_26_v_y[0+:2],_q___pip_5160_1_66___stage___block_26_v_x[0+:2]};

_t___stage___block_1280_vnum1 = {_q___pip_5160_1_66___stage___block_26_v_z[2+:2],_q___pip_5160_1_66___stage___block_26_v_y[2+:2],_q___pip_5160_1_66___stage___block_26_v_x[2+:2]};

_t___stage___block_1280_vnum2 = {_q___pip_5160_1_66___stage___block_26_v_z[4+:2],_q___pip_5160_1_66___stage___block_26_v_y[4+:2],_q___pip_5160_1_66___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_66___stage___block_6_inside&_w_tile[_t___stage___block_1280_vnum0+:1]&_w_tile[_t___stage___block_1280_vnum1+:1]&_w_tile[_t___stage___block_1280_vnum2+:1]) begin
// __block_1281
// __block_1283
_d___pip_5160_1_66___stage___block_6_clr = _t___stage___block_1280_tex;

_d___pip_5160_1_66___stage___block_6_dist = 110;

_d___pip_5160_1_66___stage___block_6_inside = 1;

// __block_1284
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1282
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1285
_t___block_1285_cmp_yx = _q___pip_5160_1_66___block_34_tm_y-_q___pip_5160_1_66___block_34_tm_x;

_t___block_1285_cmp_zx = _q___pip_5160_1_66___block_34_tm_z-_q___pip_5160_1_66___block_34_tm_x;

_t___block_1285_cmp_zy = _q___pip_5160_1_66___block_34_tm_z-_q___pip_5160_1_66___block_34_tm_y;

_t___block_1285_x_sel = ~_t___block_1285_cmp_yx[20+:1]&&~_t___block_1285_cmp_zx[20+:1];

_t___block_1285_y_sel = _t___block_1285_cmp_yx[20+:1]&&~_t___block_1285_cmp_zy[20+:1];

_t___block_1285_z_sel = _t___block_1285_cmp_zx[20+:1]&&_t___block_1285_cmp_zy[20+:1];

if (_t___block_1285_x_sel) begin
// __block_1286
// __block_1288
_d___pip_5160_1_66___stage___block_26_v_x = _q___pip_5160_1_66___stage___block_26_v_x+_q___pip_5160_1_66___stage___block_26_s_x;

_d___pip_5160_1_66___block_34_tm_x = _q___pip_5160_1_66___block_34_tm_x+_q___pip_5160_1_66___block_40_dt_x;

// __block_1289
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1287
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1290
if (_t___block_1285_y_sel) begin
// __block_1291
// __block_1293
_d___pip_5160_1_66___stage___block_26_v_y = _q___pip_5160_1_66___stage___block_26_v_y+_q___pip_5160_1_66___stage___block_26_s_y;

_d___pip_5160_1_66___block_34_tm_y = _q___pip_5160_1_66___block_34_tm_y+_q___pip_5160_1_66___block_40_dt_y;

// __block_1294
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1292
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1295
if (_t___block_1285_z_sel) begin
// __block_1296
// __block_1298
_d___pip_5160_1_66___stage___block_26_v_z = _q___pip_5160_1_66___stage___block_26_v_z+_q___pip_5160_1_66___stage___block_26_s_z;

_d___pip_5160_1_66___block_34_tm_z = _q___pip_5160_1_66___block_34_tm_z+_q___pip_5160_1_66___block_40_dt_z;

// __block_1299
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1297
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1300
// end of pipeline stage
_d__full_fsm___pip_5160_1_66 = 1;
_d__idx_fsm___pip_5160_1_66 = _t__stall_fsm___pip_5160_1_66 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_66 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 67
(* full_case *)
case (_q__idx_fsm___pip_5160_1_67)
1: begin
// __stage___block_1301
_t___stage___block_1301_tex = (_q___pip_5160_1_67___stage___block_26_v_x)^(_q___pip_5160_1_67___stage___block_26_v_y)^(_q___pip_5160_1_67___stage___block_26_v_z);

_t___stage___block_1301_vnum0 = {_q___pip_5160_1_67___stage___block_26_v_z[0+:2],_q___pip_5160_1_67___stage___block_26_v_y[0+:2],_q___pip_5160_1_67___stage___block_26_v_x[0+:2]};

_t___stage___block_1301_vnum1 = {_q___pip_5160_1_67___stage___block_26_v_z[2+:2],_q___pip_5160_1_67___stage___block_26_v_y[2+:2],_q___pip_5160_1_67___stage___block_26_v_x[2+:2]};

_t___stage___block_1301_vnum2 = {_q___pip_5160_1_67___stage___block_26_v_z[4+:2],_q___pip_5160_1_67___stage___block_26_v_y[4+:2],_q___pip_5160_1_67___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_67___stage___block_6_inside&_w_tile[_t___stage___block_1301_vnum0+:1]&_w_tile[_t___stage___block_1301_vnum1+:1]&_w_tile[_t___stage___block_1301_vnum2+:1]) begin
// __block_1302
// __block_1304
_d___pip_5160_1_67___stage___block_6_clr = _t___stage___block_1301_tex;

_d___pip_5160_1_67___stage___block_6_dist = 112;

_d___pip_5160_1_67___stage___block_6_inside = 1;

// __block_1305
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1303
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1306
_t___block_1306_cmp_yx = _q___pip_5160_1_67___block_34_tm_y-_q___pip_5160_1_67___block_34_tm_x;

_t___block_1306_cmp_zx = _q___pip_5160_1_67___block_34_tm_z-_q___pip_5160_1_67___block_34_tm_x;

_t___block_1306_cmp_zy = _q___pip_5160_1_67___block_34_tm_z-_q___pip_5160_1_67___block_34_tm_y;

_t___block_1306_x_sel = ~_t___block_1306_cmp_yx[20+:1]&&~_t___block_1306_cmp_zx[20+:1];

_t___block_1306_y_sel = _t___block_1306_cmp_yx[20+:1]&&~_t___block_1306_cmp_zy[20+:1];

_t___block_1306_z_sel = _t___block_1306_cmp_zx[20+:1]&&_t___block_1306_cmp_zy[20+:1];

if (_t___block_1306_x_sel) begin
// __block_1307
// __block_1309
_d___pip_5160_1_67___stage___block_26_v_x = _q___pip_5160_1_67___stage___block_26_v_x+_q___pip_5160_1_67___stage___block_26_s_x;

_d___pip_5160_1_67___block_34_tm_x = _q___pip_5160_1_67___block_34_tm_x+_q___pip_5160_1_67___block_40_dt_x;

// __block_1310
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1308
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1311
if (_t___block_1306_y_sel) begin
// __block_1312
// __block_1314
_d___pip_5160_1_67___stage___block_26_v_y = _q___pip_5160_1_67___stage___block_26_v_y+_q___pip_5160_1_67___stage___block_26_s_y;

_d___pip_5160_1_67___block_34_tm_y = _q___pip_5160_1_67___block_34_tm_y+_q___pip_5160_1_67___block_40_dt_y;

// __block_1315
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1313
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1316
if (_t___block_1306_z_sel) begin
// __block_1317
// __block_1319
_d___pip_5160_1_67___stage___block_26_v_z = _q___pip_5160_1_67___stage___block_26_v_z+_q___pip_5160_1_67___stage___block_26_s_z;

_d___pip_5160_1_67___block_34_tm_z = _q___pip_5160_1_67___block_34_tm_z+_q___pip_5160_1_67___block_40_dt_z;

// __block_1320
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1318
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1321
// end of pipeline stage
_d__full_fsm___pip_5160_1_67 = 1;
_d__idx_fsm___pip_5160_1_67 = _t__stall_fsm___pip_5160_1_67 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_67 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 68
(* full_case *)
case (_q__idx_fsm___pip_5160_1_68)
1: begin
// __stage___block_1322
_t___stage___block_1322_tex = (_q___pip_5160_1_68___stage___block_26_v_x)^(_q___pip_5160_1_68___stage___block_26_v_y)^(_q___pip_5160_1_68___stage___block_26_v_z);

_t___stage___block_1322_vnum0 = {_q___pip_5160_1_68___stage___block_26_v_z[0+:2],_q___pip_5160_1_68___stage___block_26_v_y[0+:2],_q___pip_5160_1_68___stage___block_26_v_x[0+:2]};

_t___stage___block_1322_vnum1 = {_q___pip_5160_1_68___stage___block_26_v_z[2+:2],_q___pip_5160_1_68___stage___block_26_v_y[2+:2],_q___pip_5160_1_68___stage___block_26_v_x[2+:2]};

_t___stage___block_1322_vnum2 = {_q___pip_5160_1_68___stage___block_26_v_z[4+:2],_q___pip_5160_1_68___stage___block_26_v_y[4+:2],_q___pip_5160_1_68___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_68___stage___block_6_inside&_w_tile[_t___stage___block_1322_vnum0+:1]&_w_tile[_t___stage___block_1322_vnum1+:1]&_w_tile[_t___stage___block_1322_vnum2+:1]) begin
// __block_1323
// __block_1325
_d___pip_5160_1_68___stage___block_6_clr = _t___stage___block_1322_tex;

_d___pip_5160_1_68___stage___block_6_dist = 113;

_d___pip_5160_1_68___stage___block_6_inside = 1;

// __block_1326
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1324
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1327
_t___block_1327_cmp_yx = _q___pip_5160_1_68___block_34_tm_y-_q___pip_5160_1_68___block_34_tm_x;

_t___block_1327_cmp_zx = _q___pip_5160_1_68___block_34_tm_z-_q___pip_5160_1_68___block_34_tm_x;

_t___block_1327_cmp_zy = _q___pip_5160_1_68___block_34_tm_z-_q___pip_5160_1_68___block_34_tm_y;

_t___block_1327_x_sel = ~_t___block_1327_cmp_yx[20+:1]&&~_t___block_1327_cmp_zx[20+:1];

_t___block_1327_y_sel = _t___block_1327_cmp_yx[20+:1]&&~_t___block_1327_cmp_zy[20+:1];

_t___block_1327_z_sel = _t___block_1327_cmp_zx[20+:1]&&_t___block_1327_cmp_zy[20+:1];

if (_t___block_1327_x_sel) begin
// __block_1328
// __block_1330
_d___pip_5160_1_68___stage___block_26_v_x = _q___pip_5160_1_68___stage___block_26_v_x+_q___pip_5160_1_68___stage___block_26_s_x;

_d___pip_5160_1_68___block_34_tm_x = _q___pip_5160_1_68___block_34_tm_x+_q___pip_5160_1_68___block_40_dt_x;

// __block_1331
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1329
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1332
if (_t___block_1327_y_sel) begin
// __block_1333
// __block_1335
_d___pip_5160_1_68___stage___block_26_v_y = _q___pip_5160_1_68___stage___block_26_v_y+_q___pip_5160_1_68___stage___block_26_s_y;

_d___pip_5160_1_68___block_34_tm_y = _q___pip_5160_1_68___block_34_tm_y+_q___pip_5160_1_68___block_40_dt_y;

// __block_1336
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1334
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1337
if (_t___block_1327_z_sel) begin
// __block_1338
// __block_1340
_d___pip_5160_1_68___stage___block_26_v_z = _q___pip_5160_1_68___stage___block_26_v_z+_q___pip_5160_1_68___stage___block_26_s_z;

_d___pip_5160_1_68___block_34_tm_z = _q___pip_5160_1_68___block_34_tm_z+_q___pip_5160_1_68___block_40_dt_z;

// __block_1341
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1339
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1342
// end of pipeline stage
_d__full_fsm___pip_5160_1_68 = 1;
_d__idx_fsm___pip_5160_1_68 = _t__stall_fsm___pip_5160_1_68 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_68 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 69
(* full_case *)
case (_q__idx_fsm___pip_5160_1_69)
1: begin
// __stage___block_1343
_t___stage___block_1343_tex = (_q___pip_5160_1_69___stage___block_26_v_x)^(_q___pip_5160_1_69___stage___block_26_v_y)^(_q___pip_5160_1_69___stage___block_26_v_z);

_t___stage___block_1343_vnum0 = {_q___pip_5160_1_69___stage___block_26_v_z[0+:2],_q___pip_5160_1_69___stage___block_26_v_y[0+:2],_q___pip_5160_1_69___stage___block_26_v_x[0+:2]};

_t___stage___block_1343_vnum1 = {_q___pip_5160_1_69___stage___block_26_v_z[2+:2],_q___pip_5160_1_69___stage___block_26_v_y[2+:2],_q___pip_5160_1_69___stage___block_26_v_x[2+:2]};

_t___stage___block_1343_vnum2 = {_q___pip_5160_1_69___stage___block_26_v_z[4+:2],_q___pip_5160_1_69___stage___block_26_v_y[4+:2],_q___pip_5160_1_69___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_69___stage___block_6_inside&_w_tile[_t___stage___block_1343_vnum0+:1]&_w_tile[_t___stage___block_1343_vnum1+:1]&_w_tile[_t___stage___block_1343_vnum2+:1]) begin
// __block_1344
// __block_1346
_d___pip_5160_1_69___stage___block_6_clr = _t___stage___block_1343_tex;

_d___pip_5160_1_69___stage___block_6_dist = 115;

_d___pip_5160_1_69___stage___block_6_inside = 1;

// __block_1347
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1345
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1348
_t___block_1348_cmp_yx = _q___pip_5160_1_69___block_34_tm_y-_q___pip_5160_1_69___block_34_tm_x;

_t___block_1348_cmp_zx = _q___pip_5160_1_69___block_34_tm_z-_q___pip_5160_1_69___block_34_tm_x;

_t___block_1348_cmp_zy = _q___pip_5160_1_69___block_34_tm_z-_q___pip_5160_1_69___block_34_tm_y;

_t___block_1348_x_sel = ~_t___block_1348_cmp_yx[20+:1]&&~_t___block_1348_cmp_zx[20+:1];

_t___block_1348_y_sel = _t___block_1348_cmp_yx[20+:1]&&~_t___block_1348_cmp_zy[20+:1];

_t___block_1348_z_sel = _t___block_1348_cmp_zx[20+:1]&&_t___block_1348_cmp_zy[20+:1];

if (_t___block_1348_x_sel) begin
// __block_1349
// __block_1351
_d___pip_5160_1_69___stage___block_26_v_x = _q___pip_5160_1_69___stage___block_26_v_x+_q___pip_5160_1_69___stage___block_26_s_x;

_d___pip_5160_1_69___block_34_tm_x = _q___pip_5160_1_69___block_34_tm_x+_q___pip_5160_1_69___block_40_dt_x;

// __block_1352
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1350
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1353
if (_t___block_1348_y_sel) begin
// __block_1354
// __block_1356
_d___pip_5160_1_69___stage___block_26_v_y = _q___pip_5160_1_69___stage___block_26_v_y+_q___pip_5160_1_69___stage___block_26_s_y;

_d___pip_5160_1_69___block_34_tm_y = _q___pip_5160_1_69___block_34_tm_y+_q___pip_5160_1_69___block_40_dt_y;

// __block_1357
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1355
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1358
if (_t___block_1348_z_sel) begin
// __block_1359
// __block_1361
_d___pip_5160_1_69___stage___block_26_v_z = _q___pip_5160_1_69___stage___block_26_v_z+_q___pip_5160_1_69___stage___block_26_s_z;

_d___pip_5160_1_69___block_34_tm_z = _q___pip_5160_1_69___block_34_tm_z+_q___pip_5160_1_69___block_40_dt_z;

// __block_1362
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1360
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1363
// end of pipeline stage
_d__full_fsm___pip_5160_1_69 = 1;
_d__idx_fsm___pip_5160_1_69 = _t__stall_fsm___pip_5160_1_69 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_69 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 70
(* full_case *)
case (_q__idx_fsm___pip_5160_1_70)
1: begin
// __stage___block_1364
_t___stage___block_1364_tex = (_q___pip_5160_1_70___stage___block_26_v_x)^(_q___pip_5160_1_70___stage___block_26_v_y)^(_q___pip_5160_1_70___stage___block_26_v_z);

_t___stage___block_1364_vnum0 = {_q___pip_5160_1_70___stage___block_26_v_z[0+:2],_q___pip_5160_1_70___stage___block_26_v_y[0+:2],_q___pip_5160_1_70___stage___block_26_v_x[0+:2]};

_t___stage___block_1364_vnum1 = {_q___pip_5160_1_70___stage___block_26_v_z[2+:2],_q___pip_5160_1_70___stage___block_26_v_y[2+:2],_q___pip_5160_1_70___stage___block_26_v_x[2+:2]};

_t___stage___block_1364_vnum2 = {_q___pip_5160_1_70___stage___block_26_v_z[4+:2],_q___pip_5160_1_70___stage___block_26_v_y[4+:2],_q___pip_5160_1_70___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_70___stage___block_6_inside&_w_tile[_t___stage___block_1364_vnum0+:1]&_w_tile[_t___stage___block_1364_vnum1+:1]&_w_tile[_t___stage___block_1364_vnum2+:1]) begin
// __block_1365
// __block_1367
_d___pip_5160_1_70___stage___block_6_clr = _t___stage___block_1364_tex;

_d___pip_5160_1_70___stage___block_6_dist = 117;

_d___pip_5160_1_70___stage___block_6_inside = 1;

// __block_1368
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1366
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1369
_t___block_1369_cmp_yx = _q___pip_5160_1_70___block_34_tm_y-_q___pip_5160_1_70___block_34_tm_x;

_t___block_1369_cmp_zx = _q___pip_5160_1_70___block_34_tm_z-_q___pip_5160_1_70___block_34_tm_x;

_t___block_1369_cmp_zy = _q___pip_5160_1_70___block_34_tm_z-_q___pip_5160_1_70___block_34_tm_y;

_t___block_1369_x_sel = ~_t___block_1369_cmp_yx[20+:1]&&~_t___block_1369_cmp_zx[20+:1];

_t___block_1369_y_sel = _t___block_1369_cmp_yx[20+:1]&&~_t___block_1369_cmp_zy[20+:1];

_t___block_1369_z_sel = _t___block_1369_cmp_zx[20+:1]&&_t___block_1369_cmp_zy[20+:1];

if (_t___block_1369_x_sel) begin
// __block_1370
// __block_1372
_d___pip_5160_1_70___stage___block_26_v_x = _q___pip_5160_1_70___stage___block_26_v_x+_q___pip_5160_1_70___stage___block_26_s_x;

_d___pip_5160_1_70___block_34_tm_x = _q___pip_5160_1_70___block_34_tm_x+_q___pip_5160_1_70___block_40_dt_x;

// __block_1373
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1371
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1374
if (_t___block_1369_y_sel) begin
// __block_1375
// __block_1377
_d___pip_5160_1_70___stage___block_26_v_y = _q___pip_5160_1_70___stage___block_26_v_y+_q___pip_5160_1_70___stage___block_26_s_y;

_d___pip_5160_1_70___block_34_tm_y = _q___pip_5160_1_70___block_34_tm_y+_q___pip_5160_1_70___block_40_dt_y;

// __block_1378
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1376
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1379
if (_t___block_1369_z_sel) begin
// __block_1380
// __block_1382
_d___pip_5160_1_70___stage___block_26_v_z = _q___pip_5160_1_70___stage___block_26_v_z+_q___pip_5160_1_70___stage___block_26_s_z;

_d___pip_5160_1_70___block_34_tm_z = _q___pip_5160_1_70___block_34_tm_z+_q___pip_5160_1_70___block_40_dt_z;

// __block_1383
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1381
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1384
// end of pipeline stage
_d__full_fsm___pip_5160_1_70 = 1;
_d__idx_fsm___pip_5160_1_70 = _t__stall_fsm___pip_5160_1_70 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_70 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 71
(* full_case *)
case (_q__idx_fsm___pip_5160_1_71)
1: begin
// __stage___block_1385
_t___stage___block_1385_tex = (_q___pip_5160_1_71___stage___block_26_v_x)^(_q___pip_5160_1_71___stage___block_26_v_y)^(_q___pip_5160_1_71___stage___block_26_v_z);

_t___stage___block_1385_vnum0 = {_q___pip_5160_1_71___stage___block_26_v_z[0+:2],_q___pip_5160_1_71___stage___block_26_v_y[0+:2],_q___pip_5160_1_71___stage___block_26_v_x[0+:2]};

_t___stage___block_1385_vnum1 = {_q___pip_5160_1_71___stage___block_26_v_z[2+:2],_q___pip_5160_1_71___stage___block_26_v_y[2+:2],_q___pip_5160_1_71___stage___block_26_v_x[2+:2]};

_t___stage___block_1385_vnum2 = {_q___pip_5160_1_71___stage___block_26_v_z[4+:2],_q___pip_5160_1_71___stage___block_26_v_y[4+:2],_q___pip_5160_1_71___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_71___stage___block_6_inside&_w_tile[_t___stage___block_1385_vnum0+:1]&_w_tile[_t___stage___block_1385_vnum1+:1]&_w_tile[_t___stage___block_1385_vnum2+:1]) begin
// __block_1386
// __block_1388
_d___pip_5160_1_71___stage___block_6_clr = _t___stage___block_1385_tex;

_d___pip_5160_1_71___stage___block_6_dist = 119;

_d___pip_5160_1_71___stage___block_6_inside = 1;

// __block_1389
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1387
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1390
_t___block_1390_cmp_yx = _q___pip_5160_1_71___block_34_tm_y-_q___pip_5160_1_71___block_34_tm_x;

_t___block_1390_cmp_zx = _q___pip_5160_1_71___block_34_tm_z-_q___pip_5160_1_71___block_34_tm_x;

_t___block_1390_cmp_zy = _q___pip_5160_1_71___block_34_tm_z-_q___pip_5160_1_71___block_34_tm_y;

_t___block_1390_x_sel = ~_t___block_1390_cmp_yx[20+:1]&&~_t___block_1390_cmp_zx[20+:1];

_t___block_1390_y_sel = _t___block_1390_cmp_yx[20+:1]&&~_t___block_1390_cmp_zy[20+:1];

_t___block_1390_z_sel = _t___block_1390_cmp_zx[20+:1]&&_t___block_1390_cmp_zy[20+:1];

if (_t___block_1390_x_sel) begin
// __block_1391
// __block_1393
_d___pip_5160_1_71___stage___block_26_v_x = _q___pip_5160_1_71___stage___block_26_v_x+_q___pip_5160_1_71___stage___block_26_s_x;

_d___pip_5160_1_71___block_34_tm_x = _q___pip_5160_1_71___block_34_tm_x+_q___pip_5160_1_71___block_40_dt_x;

// __block_1394
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1392
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1395
if (_t___block_1390_y_sel) begin
// __block_1396
// __block_1398
_d___pip_5160_1_71___stage___block_26_v_y = _q___pip_5160_1_71___stage___block_26_v_y+_q___pip_5160_1_71___stage___block_26_s_y;

_d___pip_5160_1_71___block_34_tm_y = _q___pip_5160_1_71___block_34_tm_y+_q___pip_5160_1_71___block_40_dt_y;

// __block_1399
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1397
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1400
if (_t___block_1390_z_sel) begin
// __block_1401
// __block_1403
_d___pip_5160_1_71___stage___block_26_v_z = _q___pip_5160_1_71___stage___block_26_v_z+_q___pip_5160_1_71___stage___block_26_s_z;

_d___pip_5160_1_71___block_34_tm_z = _q___pip_5160_1_71___block_34_tm_z+_q___pip_5160_1_71___block_40_dt_z;

// __block_1404
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1402
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1405
// end of pipeline stage
_d__full_fsm___pip_5160_1_71 = 1;
_d__idx_fsm___pip_5160_1_71 = _t__stall_fsm___pip_5160_1_71 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_71 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 72
(* full_case *)
case (_q__idx_fsm___pip_5160_1_72)
1: begin
// __stage___block_1406
_t___stage___block_1406_tex = (_q___pip_5160_1_72___stage___block_26_v_x)^(_q___pip_5160_1_72___stage___block_26_v_y)^(_q___pip_5160_1_72___stage___block_26_v_z);

_t___stage___block_1406_vnum0 = {_q___pip_5160_1_72___stage___block_26_v_z[0+:2],_q___pip_5160_1_72___stage___block_26_v_y[0+:2],_q___pip_5160_1_72___stage___block_26_v_x[0+:2]};

_t___stage___block_1406_vnum1 = {_q___pip_5160_1_72___stage___block_26_v_z[2+:2],_q___pip_5160_1_72___stage___block_26_v_y[2+:2],_q___pip_5160_1_72___stage___block_26_v_x[2+:2]};

_t___stage___block_1406_vnum2 = {_q___pip_5160_1_72___stage___block_26_v_z[4+:2],_q___pip_5160_1_72___stage___block_26_v_y[4+:2],_q___pip_5160_1_72___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_72___stage___block_6_inside&_w_tile[_t___stage___block_1406_vnum0+:1]&_w_tile[_t___stage___block_1406_vnum1+:1]&_w_tile[_t___stage___block_1406_vnum2+:1]) begin
// __block_1407
// __block_1409
_d___pip_5160_1_72___stage___block_6_clr = _t___stage___block_1406_tex;

_d___pip_5160_1_72___stage___block_6_dist = 121;

_d___pip_5160_1_72___stage___block_6_inside = 1;

// __block_1410
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1408
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1411
_t___block_1411_cmp_yx = _q___pip_5160_1_72___block_34_tm_y-_q___pip_5160_1_72___block_34_tm_x;

_t___block_1411_cmp_zx = _q___pip_5160_1_72___block_34_tm_z-_q___pip_5160_1_72___block_34_tm_x;

_t___block_1411_cmp_zy = _q___pip_5160_1_72___block_34_tm_z-_q___pip_5160_1_72___block_34_tm_y;

_t___block_1411_x_sel = ~_t___block_1411_cmp_yx[20+:1]&&~_t___block_1411_cmp_zx[20+:1];

_t___block_1411_y_sel = _t___block_1411_cmp_yx[20+:1]&&~_t___block_1411_cmp_zy[20+:1];

_t___block_1411_z_sel = _t___block_1411_cmp_zx[20+:1]&&_t___block_1411_cmp_zy[20+:1];

if (_t___block_1411_x_sel) begin
// __block_1412
// __block_1414
_d___pip_5160_1_72___stage___block_26_v_x = _q___pip_5160_1_72___stage___block_26_v_x+_q___pip_5160_1_72___stage___block_26_s_x;

_d___pip_5160_1_72___block_34_tm_x = _q___pip_5160_1_72___block_34_tm_x+_q___pip_5160_1_72___block_40_dt_x;

// __block_1415
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1413
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1416
if (_t___block_1411_y_sel) begin
// __block_1417
// __block_1419
_d___pip_5160_1_72___stage___block_26_v_y = _q___pip_5160_1_72___stage___block_26_v_y+_q___pip_5160_1_72___stage___block_26_s_y;

_d___pip_5160_1_72___block_34_tm_y = _q___pip_5160_1_72___block_34_tm_y+_q___pip_5160_1_72___block_40_dt_y;

// __block_1420
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1418
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1421
if (_t___block_1411_z_sel) begin
// __block_1422
// __block_1424
_d___pip_5160_1_72___stage___block_26_v_z = _q___pip_5160_1_72___stage___block_26_v_z+_q___pip_5160_1_72___stage___block_26_s_z;

_d___pip_5160_1_72___block_34_tm_z = _q___pip_5160_1_72___block_34_tm_z+_q___pip_5160_1_72___block_40_dt_z;

// __block_1425
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1423
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1426
// end of pipeline stage
_d__full_fsm___pip_5160_1_72 = 1;
_d__idx_fsm___pip_5160_1_72 = _t__stall_fsm___pip_5160_1_72 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_72 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 73
(* full_case *)
case (_q__idx_fsm___pip_5160_1_73)
1: begin
// __stage___block_1427
_t___stage___block_1427_tex = (_q___pip_5160_1_73___stage___block_26_v_x)^(_q___pip_5160_1_73___stage___block_26_v_y)^(_q___pip_5160_1_73___stage___block_26_v_z);

_t___stage___block_1427_vnum0 = {_q___pip_5160_1_73___stage___block_26_v_z[0+:2],_q___pip_5160_1_73___stage___block_26_v_y[0+:2],_q___pip_5160_1_73___stage___block_26_v_x[0+:2]};

_t___stage___block_1427_vnum1 = {_q___pip_5160_1_73___stage___block_26_v_z[2+:2],_q___pip_5160_1_73___stage___block_26_v_y[2+:2],_q___pip_5160_1_73___stage___block_26_v_x[2+:2]};

_t___stage___block_1427_vnum2 = {_q___pip_5160_1_73___stage___block_26_v_z[4+:2],_q___pip_5160_1_73___stage___block_26_v_y[4+:2],_q___pip_5160_1_73___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_73___stage___block_6_inside&_w_tile[_t___stage___block_1427_vnum0+:1]&_w_tile[_t___stage___block_1427_vnum1+:1]&_w_tile[_t___stage___block_1427_vnum2+:1]) begin
// __block_1428
// __block_1430
_d___pip_5160_1_73___stage___block_6_clr = _t___stage___block_1427_tex;

_d___pip_5160_1_73___stage___block_6_dist = 123;

_d___pip_5160_1_73___stage___block_6_inside = 1;

// __block_1431
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1429
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1432
_t___block_1432_cmp_yx = _q___pip_5160_1_73___block_34_tm_y-_q___pip_5160_1_73___block_34_tm_x;

_t___block_1432_cmp_zx = _q___pip_5160_1_73___block_34_tm_z-_q___pip_5160_1_73___block_34_tm_x;

_t___block_1432_cmp_zy = _q___pip_5160_1_73___block_34_tm_z-_q___pip_5160_1_73___block_34_tm_y;

_t___block_1432_x_sel = ~_t___block_1432_cmp_yx[20+:1]&&~_t___block_1432_cmp_zx[20+:1];

_t___block_1432_y_sel = _t___block_1432_cmp_yx[20+:1]&&~_t___block_1432_cmp_zy[20+:1];

_t___block_1432_z_sel = _t___block_1432_cmp_zx[20+:1]&&_t___block_1432_cmp_zy[20+:1];

if (_t___block_1432_x_sel) begin
// __block_1433
// __block_1435
_d___pip_5160_1_73___stage___block_26_v_x = _q___pip_5160_1_73___stage___block_26_v_x+_q___pip_5160_1_73___stage___block_26_s_x;

_d___pip_5160_1_73___block_34_tm_x = _q___pip_5160_1_73___block_34_tm_x+_q___pip_5160_1_73___block_40_dt_x;

// __block_1436
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1434
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1437
if (_t___block_1432_y_sel) begin
// __block_1438
// __block_1440
_d___pip_5160_1_73___stage___block_26_v_y = _q___pip_5160_1_73___stage___block_26_v_y+_q___pip_5160_1_73___stage___block_26_s_y;

_d___pip_5160_1_73___block_34_tm_y = _q___pip_5160_1_73___block_34_tm_y+_q___pip_5160_1_73___block_40_dt_y;

// __block_1441
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1439
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1442
if (_t___block_1432_z_sel) begin
// __block_1443
// __block_1445
_d___pip_5160_1_73___stage___block_26_v_z = _q___pip_5160_1_73___stage___block_26_v_z+_q___pip_5160_1_73___stage___block_26_s_z;

_d___pip_5160_1_73___block_34_tm_z = _q___pip_5160_1_73___block_34_tm_z+_q___pip_5160_1_73___block_40_dt_z;

// __block_1446
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1444
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1447
// end of pipeline stage
_d__full_fsm___pip_5160_1_73 = 1;
_d__idx_fsm___pip_5160_1_73 = _t__stall_fsm___pip_5160_1_73 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_73 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 74
(* full_case *)
case (_q__idx_fsm___pip_5160_1_74)
1: begin
// __stage___block_1448
_t___stage___block_1448_tex = (_q___pip_5160_1_74___stage___block_26_v_x)^(_q___pip_5160_1_74___stage___block_26_v_y)^(_q___pip_5160_1_74___stage___block_26_v_z);

_t___stage___block_1448_vnum0 = {_q___pip_5160_1_74___stage___block_26_v_z[0+:2],_q___pip_5160_1_74___stage___block_26_v_y[0+:2],_q___pip_5160_1_74___stage___block_26_v_x[0+:2]};

_t___stage___block_1448_vnum1 = {_q___pip_5160_1_74___stage___block_26_v_z[2+:2],_q___pip_5160_1_74___stage___block_26_v_y[2+:2],_q___pip_5160_1_74___stage___block_26_v_x[2+:2]};

_t___stage___block_1448_vnum2 = {_q___pip_5160_1_74___stage___block_26_v_z[4+:2],_q___pip_5160_1_74___stage___block_26_v_y[4+:2],_q___pip_5160_1_74___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_74___stage___block_6_inside&_w_tile[_t___stage___block_1448_vnum0+:1]&_w_tile[_t___stage___block_1448_vnum1+:1]&_w_tile[_t___stage___block_1448_vnum2+:1]) begin
// __block_1449
// __block_1451
_d___pip_5160_1_74___stage___block_6_clr = _t___stage___block_1448_tex;

_d___pip_5160_1_74___stage___block_6_dist = 125;

_d___pip_5160_1_74___stage___block_6_inside = 1;

// __block_1452
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1450
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1453
_t___block_1453_cmp_yx = _q___pip_5160_1_74___block_34_tm_y-_q___pip_5160_1_74___block_34_tm_x;

_t___block_1453_cmp_zx = _q___pip_5160_1_74___block_34_tm_z-_q___pip_5160_1_74___block_34_tm_x;

_t___block_1453_cmp_zy = _q___pip_5160_1_74___block_34_tm_z-_q___pip_5160_1_74___block_34_tm_y;

_t___block_1453_x_sel = ~_t___block_1453_cmp_yx[20+:1]&&~_t___block_1453_cmp_zx[20+:1];

_t___block_1453_y_sel = _t___block_1453_cmp_yx[20+:1]&&~_t___block_1453_cmp_zy[20+:1];

_t___block_1453_z_sel = _t___block_1453_cmp_zx[20+:1]&&_t___block_1453_cmp_zy[20+:1];

if (_t___block_1453_x_sel) begin
// __block_1454
// __block_1456
_d___pip_5160_1_74___stage___block_26_v_x = _q___pip_5160_1_74___stage___block_26_v_x+_q___pip_5160_1_74___stage___block_26_s_x;

_d___pip_5160_1_74___block_34_tm_x = _q___pip_5160_1_74___block_34_tm_x+_q___pip_5160_1_74___block_40_dt_x;

// __block_1457
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1455
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1458
if (_t___block_1453_y_sel) begin
// __block_1459
// __block_1461
_d___pip_5160_1_74___stage___block_26_v_y = _q___pip_5160_1_74___stage___block_26_v_y+_q___pip_5160_1_74___stage___block_26_s_y;

_d___pip_5160_1_74___block_34_tm_y = _q___pip_5160_1_74___block_34_tm_y+_q___pip_5160_1_74___block_40_dt_y;

// __block_1462
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1460
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1463
if (_t___block_1453_z_sel) begin
// __block_1464
// __block_1466
_d___pip_5160_1_74___stage___block_26_v_z = _q___pip_5160_1_74___stage___block_26_v_z+_q___pip_5160_1_74___stage___block_26_s_z;

_d___pip_5160_1_74___block_34_tm_z = _q___pip_5160_1_74___block_34_tm_z+_q___pip_5160_1_74___block_40_dt_z;

// __block_1467
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1465
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1468
// end of pipeline stage
_d__full_fsm___pip_5160_1_74 = 1;
_d__idx_fsm___pip_5160_1_74 = _t__stall_fsm___pip_5160_1_74 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_74 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 75
(* full_case *)
case (_q__idx_fsm___pip_5160_1_75)
1: begin
// __stage___block_1469
_t___stage___block_1469_tex = (_q___pip_5160_1_75___stage___block_26_v_x)^(_q___pip_5160_1_75___stage___block_26_v_y)^(_q___pip_5160_1_75___stage___block_26_v_z);

_t___stage___block_1469_vnum0 = {_q___pip_5160_1_75___stage___block_26_v_z[0+:2],_q___pip_5160_1_75___stage___block_26_v_y[0+:2],_q___pip_5160_1_75___stage___block_26_v_x[0+:2]};

_t___stage___block_1469_vnum1 = {_q___pip_5160_1_75___stage___block_26_v_z[2+:2],_q___pip_5160_1_75___stage___block_26_v_y[2+:2],_q___pip_5160_1_75___stage___block_26_v_x[2+:2]};

_t___stage___block_1469_vnum2 = {_q___pip_5160_1_75___stage___block_26_v_z[4+:2],_q___pip_5160_1_75___stage___block_26_v_y[4+:2],_q___pip_5160_1_75___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_75___stage___block_6_inside&_w_tile[_t___stage___block_1469_vnum0+:1]&_w_tile[_t___stage___block_1469_vnum1+:1]&_w_tile[_t___stage___block_1469_vnum2+:1]) begin
// __block_1470
// __block_1472
_d___pip_5160_1_75___stage___block_6_clr = _t___stage___block_1469_tex;

_d___pip_5160_1_75___stage___block_6_dist = 126;

_d___pip_5160_1_75___stage___block_6_inside = 1;

// __block_1473
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1471
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1474
_t___block_1474_cmp_yx = _q___pip_5160_1_75___block_34_tm_y-_q___pip_5160_1_75___block_34_tm_x;

_t___block_1474_cmp_zx = _q___pip_5160_1_75___block_34_tm_z-_q___pip_5160_1_75___block_34_tm_x;

_t___block_1474_cmp_zy = _q___pip_5160_1_75___block_34_tm_z-_q___pip_5160_1_75___block_34_tm_y;

_t___block_1474_x_sel = ~_t___block_1474_cmp_yx[20+:1]&&~_t___block_1474_cmp_zx[20+:1];

_t___block_1474_y_sel = _t___block_1474_cmp_yx[20+:1]&&~_t___block_1474_cmp_zy[20+:1];

_t___block_1474_z_sel = _t___block_1474_cmp_zx[20+:1]&&_t___block_1474_cmp_zy[20+:1];

if (_t___block_1474_x_sel) begin
// __block_1475
// __block_1477
_d___pip_5160_1_75___stage___block_26_v_x = _q___pip_5160_1_75___stage___block_26_v_x+_q___pip_5160_1_75___stage___block_26_s_x;

_d___pip_5160_1_75___block_34_tm_x = _q___pip_5160_1_75___block_34_tm_x+_q___pip_5160_1_75___block_40_dt_x;

// __block_1478
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1476
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1479
if (_t___block_1474_y_sel) begin
// __block_1480
// __block_1482
_d___pip_5160_1_75___stage___block_26_v_y = _q___pip_5160_1_75___stage___block_26_v_y+_q___pip_5160_1_75___stage___block_26_s_y;

_d___pip_5160_1_75___block_34_tm_y = _q___pip_5160_1_75___block_34_tm_y+_q___pip_5160_1_75___block_40_dt_y;

// __block_1483
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1481
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1484
if (_t___block_1474_z_sel) begin
// __block_1485
// __block_1487
_d___pip_5160_1_75___stage___block_26_v_z = _q___pip_5160_1_75___stage___block_26_v_z+_q___pip_5160_1_75___stage___block_26_s_z;

_d___pip_5160_1_75___block_34_tm_z = _q___pip_5160_1_75___block_34_tm_z+_q___pip_5160_1_75___block_40_dt_z;

// __block_1488
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1486
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1489
// end of pipeline stage
_d__full_fsm___pip_5160_1_75 = 1;
_d__idx_fsm___pip_5160_1_75 = _t__stall_fsm___pip_5160_1_75 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_75 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 76
(* full_case *)
case (_q__idx_fsm___pip_5160_1_76)
1: begin
// __stage___block_1490
_t___stage___block_1490_tex = (_q___pip_5160_1_76___stage___block_26_v_x)^(_q___pip_5160_1_76___stage___block_26_v_y)^(_q___pip_5160_1_76___stage___block_26_v_z);

_t___stage___block_1490_vnum0 = {_q___pip_5160_1_76___stage___block_26_v_z[0+:2],_q___pip_5160_1_76___stage___block_26_v_y[0+:2],_q___pip_5160_1_76___stage___block_26_v_x[0+:2]};

_t___stage___block_1490_vnum1 = {_q___pip_5160_1_76___stage___block_26_v_z[2+:2],_q___pip_5160_1_76___stage___block_26_v_y[2+:2],_q___pip_5160_1_76___stage___block_26_v_x[2+:2]};

_t___stage___block_1490_vnum2 = {_q___pip_5160_1_76___stage___block_26_v_z[4+:2],_q___pip_5160_1_76___stage___block_26_v_y[4+:2],_q___pip_5160_1_76___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_76___stage___block_6_inside&_w_tile[_t___stage___block_1490_vnum0+:1]&_w_tile[_t___stage___block_1490_vnum1+:1]&_w_tile[_t___stage___block_1490_vnum2+:1]) begin
// __block_1491
// __block_1493
_d___pip_5160_1_76___stage___block_6_clr = _t___stage___block_1490_tex;

_d___pip_5160_1_76___stage___block_6_dist = 128;

_d___pip_5160_1_76___stage___block_6_inside = 1;

// __block_1494
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1492
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1495
_t___block_1495_cmp_yx = _q___pip_5160_1_76___block_34_tm_y-_q___pip_5160_1_76___block_34_tm_x;

_t___block_1495_cmp_zx = _q___pip_5160_1_76___block_34_tm_z-_q___pip_5160_1_76___block_34_tm_x;

_t___block_1495_cmp_zy = _q___pip_5160_1_76___block_34_tm_z-_q___pip_5160_1_76___block_34_tm_y;

_t___block_1495_x_sel = ~_t___block_1495_cmp_yx[20+:1]&&~_t___block_1495_cmp_zx[20+:1];

_t___block_1495_y_sel = _t___block_1495_cmp_yx[20+:1]&&~_t___block_1495_cmp_zy[20+:1];

_t___block_1495_z_sel = _t___block_1495_cmp_zx[20+:1]&&_t___block_1495_cmp_zy[20+:1];

if (_t___block_1495_x_sel) begin
// __block_1496
// __block_1498
_d___pip_5160_1_76___stage___block_26_v_x = _q___pip_5160_1_76___stage___block_26_v_x+_q___pip_5160_1_76___stage___block_26_s_x;

_d___pip_5160_1_76___block_34_tm_x = _q___pip_5160_1_76___block_34_tm_x+_q___pip_5160_1_76___block_40_dt_x;

// __block_1499
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1497
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1500
if (_t___block_1495_y_sel) begin
// __block_1501
// __block_1503
_d___pip_5160_1_76___stage___block_26_v_y = _q___pip_5160_1_76___stage___block_26_v_y+_q___pip_5160_1_76___stage___block_26_s_y;

_d___pip_5160_1_76___block_34_tm_y = _q___pip_5160_1_76___block_34_tm_y+_q___pip_5160_1_76___block_40_dt_y;

// __block_1504
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1502
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1505
if (_t___block_1495_z_sel) begin
// __block_1506
// __block_1508
_d___pip_5160_1_76___stage___block_26_v_z = _q___pip_5160_1_76___stage___block_26_v_z+_q___pip_5160_1_76___stage___block_26_s_z;

_d___pip_5160_1_76___block_34_tm_z = _q___pip_5160_1_76___block_34_tm_z+_q___pip_5160_1_76___block_40_dt_z;

// __block_1509
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1507
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1510
// end of pipeline stage
_d__full_fsm___pip_5160_1_76 = 1;
_d__idx_fsm___pip_5160_1_76 = _t__stall_fsm___pip_5160_1_76 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_76 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 77
(* full_case *)
case (_q__idx_fsm___pip_5160_1_77)
1: begin
// __stage___block_1511
_t___stage___block_1511_tex = (_q___pip_5160_1_77___stage___block_26_v_x)^(_q___pip_5160_1_77___stage___block_26_v_y)^(_q___pip_5160_1_77___stage___block_26_v_z);

_t___stage___block_1511_vnum0 = {_q___pip_5160_1_77___stage___block_26_v_z[0+:2],_q___pip_5160_1_77___stage___block_26_v_y[0+:2],_q___pip_5160_1_77___stage___block_26_v_x[0+:2]};

_t___stage___block_1511_vnum1 = {_q___pip_5160_1_77___stage___block_26_v_z[2+:2],_q___pip_5160_1_77___stage___block_26_v_y[2+:2],_q___pip_5160_1_77___stage___block_26_v_x[2+:2]};

_t___stage___block_1511_vnum2 = {_q___pip_5160_1_77___stage___block_26_v_z[4+:2],_q___pip_5160_1_77___stage___block_26_v_y[4+:2],_q___pip_5160_1_77___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_77___stage___block_6_inside&_w_tile[_t___stage___block_1511_vnum0+:1]&_w_tile[_t___stage___block_1511_vnum1+:1]&_w_tile[_t___stage___block_1511_vnum2+:1]) begin
// __block_1512
// __block_1514
_d___pip_5160_1_77___stage___block_6_clr = _t___stage___block_1511_tex;

_d___pip_5160_1_77___stage___block_6_dist = 130;

_d___pip_5160_1_77___stage___block_6_inside = 1;

// __block_1515
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1513
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1516
_t___block_1516_cmp_yx = _q___pip_5160_1_77___block_34_tm_y-_q___pip_5160_1_77___block_34_tm_x;

_t___block_1516_cmp_zx = _q___pip_5160_1_77___block_34_tm_z-_q___pip_5160_1_77___block_34_tm_x;

_t___block_1516_cmp_zy = _q___pip_5160_1_77___block_34_tm_z-_q___pip_5160_1_77___block_34_tm_y;

_t___block_1516_x_sel = ~_t___block_1516_cmp_yx[20+:1]&&~_t___block_1516_cmp_zx[20+:1];

_t___block_1516_y_sel = _t___block_1516_cmp_yx[20+:1]&&~_t___block_1516_cmp_zy[20+:1];

_t___block_1516_z_sel = _t___block_1516_cmp_zx[20+:1]&&_t___block_1516_cmp_zy[20+:1];

if (_t___block_1516_x_sel) begin
// __block_1517
// __block_1519
_d___pip_5160_1_77___stage___block_26_v_x = _q___pip_5160_1_77___stage___block_26_v_x+_q___pip_5160_1_77___stage___block_26_s_x;

_d___pip_5160_1_77___block_34_tm_x = _q___pip_5160_1_77___block_34_tm_x+_q___pip_5160_1_77___block_40_dt_x;

// __block_1520
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1518
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1521
if (_t___block_1516_y_sel) begin
// __block_1522
// __block_1524
_d___pip_5160_1_77___stage___block_26_v_y = _q___pip_5160_1_77___stage___block_26_v_y+_q___pip_5160_1_77___stage___block_26_s_y;

_d___pip_5160_1_77___block_34_tm_y = _q___pip_5160_1_77___block_34_tm_y+_q___pip_5160_1_77___block_40_dt_y;

// __block_1525
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1523
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1526
if (_t___block_1516_z_sel) begin
// __block_1527
// __block_1529
_d___pip_5160_1_77___stage___block_26_v_z = _q___pip_5160_1_77___stage___block_26_v_z+_q___pip_5160_1_77___stage___block_26_s_z;

_d___pip_5160_1_77___block_34_tm_z = _q___pip_5160_1_77___block_34_tm_z+_q___pip_5160_1_77___block_40_dt_z;

// __block_1530
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1528
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1531
// end of pipeline stage
_d__full_fsm___pip_5160_1_77 = 1;
_d__idx_fsm___pip_5160_1_77 = _t__stall_fsm___pip_5160_1_77 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_77 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 78
(* full_case *)
case (_q__idx_fsm___pip_5160_1_78)
1: begin
// __stage___block_1532
_t___stage___block_1532_tex = (_q___pip_5160_1_78___stage___block_26_v_x)^(_q___pip_5160_1_78___stage___block_26_v_y)^(_q___pip_5160_1_78___stage___block_26_v_z);

_t___stage___block_1532_vnum0 = {_q___pip_5160_1_78___stage___block_26_v_z[0+:2],_q___pip_5160_1_78___stage___block_26_v_y[0+:2],_q___pip_5160_1_78___stage___block_26_v_x[0+:2]};

_t___stage___block_1532_vnum1 = {_q___pip_5160_1_78___stage___block_26_v_z[2+:2],_q___pip_5160_1_78___stage___block_26_v_y[2+:2],_q___pip_5160_1_78___stage___block_26_v_x[2+:2]};

_t___stage___block_1532_vnum2 = {_q___pip_5160_1_78___stage___block_26_v_z[4+:2],_q___pip_5160_1_78___stage___block_26_v_y[4+:2],_q___pip_5160_1_78___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_78___stage___block_6_inside&_w_tile[_t___stage___block_1532_vnum0+:1]&_w_tile[_t___stage___block_1532_vnum1+:1]&_w_tile[_t___stage___block_1532_vnum2+:1]) begin
// __block_1533
// __block_1535
_d___pip_5160_1_78___stage___block_6_clr = _t___stage___block_1532_tex;

_d___pip_5160_1_78___stage___block_6_dist = 132;

_d___pip_5160_1_78___stage___block_6_inside = 1;

// __block_1536
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1534
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1537
_t___block_1537_cmp_yx = _q___pip_5160_1_78___block_34_tm_y-_q___pip_5160_1_78___block_34_tm_x;

_t___block_1537_cmp_zx = _q___pip_5160_1_78___block_34_tm_z-_q___pip_5160_1_78___block_34_tm_x;

_t___block_1537_cmp_zy = _q___pip_5160_1_78___block_34_tm_z-_q___pip_5160_1_78___block_34_tm_y;

_t___block_1537_x_sel = ~_t___block_1537_cmp_yx[20+:1]&&~_t___block_1537_cmp_zx[20+:1];

_t___block_1537_y_sel = _t___block_1537_cmp_yx[20+:1]&&~_t___block_1537_cmp_zy[20+:1];

_t___block_1537_z_sel = _t___block_1537_cmp_zx[20+:1]&&_t___block_1537_cmp_zy[20+:1];

if (_t___block_1537_x_sel) begin
// __block_1538
// __block_1540
_d___pip_5160_1_78___stage___block_26_v_x = _q___pip_5160_1_78___stage___block_26_v_x+_q___pip_5160_1_78___stage___block_26_s_x;

_d___pip_5160_1_78___block_34_tm_x = _q___pip_5160_1_78___block_34_tm_x+_q___pip_5160_1_78___block_40_dt_x;

// __block_1541
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1539
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1542
if (_t___block_1537_y_sel) begin
// __block_1543
// __block_1545
_d___pip_5160_1_78___stage___block_26_v_y = _q___pip_5160_1_78___stage___block_26_v_y+_q___pip_5160_1_78___stage___block_26_s_y;

_d___pip_5160_1_78___block_34_tm_y = _q___pip_5160_1_78___block_34_tm_y+_q___pip_5160_1_78___block_40_dt_y;

// __block_1546
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1544
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1547
if (_t___block_1537_z_sel) begin
// __block_1548
// __block_1550
_d___pip_5160_1_78___stage___block_26_v_z = _q___pip_5160_1_78___stage___block_26_v_z+_q___pip_5160_1_78___stage___block_26_s_z;

_d___pip_5160_1_78___block_34_tm_z = _q___pip_5160_1_78___block_34_tm_z+_q___pip_5160_1_78___block_40_dt_z;

// __block_1551
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1549
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1552
// end of pipeline stage
_d__full_fsm___pip_5160_1_78 = 1;
_d__idx_fsm___pip_5160_1_78 = _t__stall_fsm___pip_5160_1_78 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_78 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 79
(* full_case *)
case (_q__idx_fsm___pip_5160_1_79)
1: begin
// __stage___block_1553
_t___stage___block_1553_tex = (_q___pip_5160_1_79___stage___block_26_v_x)^(_q___pip_5160_1_79___stage___block_26_v_y)^(_q___pip_5160_1_79___stage___block_26_v_z);

_t___stage___block_1553_vnum0 = {_q___pip_5160_1_79___stage___block_26_v_z[0+:2],_q___pip_5160_1_79___stage___block_26_v_y[0+:2],_q___pip_5160_1_79___stage___block_26_v_x[0+:2]};

_t___stage___block_1553_vnum1 = {_q___pip_5160_1_79___stage___block_26_v_z[2+:2],_q___pip_5160_1_79___stage___block_26_v_y[2+:2],_q___pip_5160_1_79___stage___block_26_v_x[2+:2]};

_t___stage___block_1553_vnum2 = {_q___pip_5160_1_79___stage___block_26_v_z[4+:2],_q___pip_5160_1_79___stage___block_26_v_y[4+:2],_q___pip_5160_1_79___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_79___stage___block_6_inside&_w_tile[_t___stage___block_1553_vnum0+:1]&_w_tile[_t___stage___block_1553_vnum1+:1]&_w_tile[_t___stage___block_1553_vnum2+:1]) begin
// __block_1554
// __block_1556
_d___pip_5160_1_79___stage___block_6_clr = _t___stage___block_1553_tex;

_d___pip_5160_1_79___stage___block_6_dist = 134;

_d___pip_5160_1_79___stage___block_6_inside = 1;

// __block_1557
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1555
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1558
_t___block_1558_cmp_yx = _q___pip_5160_1_79___block_34_tm_y-_q___pip_5160_1_79___block_34_tm_x;

_t___block_1558_cmp_zx = _q___pip_5160_1_79___block_34_tm_z-_q___pip_5160_1_79___block_34_tm_x;

_t___block_1558_cmp_zy = _q___pip_5160_1_79___block_34_tm_z-_q___pip_5160_1_79___block_34_tm_y;

_t___block_1558_x_sel = ~_t___block_1558_cmp_yx[20+:1]&&~_t___block_1558_cmp_zx[20+:1];

_t___block_1558_y_sel = _t___block_1558_cmp_yx[20+:1]&&~_t___block_1558_cmp_zy[20+:1];

_t___block_1558_z_sel = _t___block_1558_cmp_zx[20+:1]&&_t___block_1558_cmp_zy[20+:1];

if (_t___block_1558_x_sel) begin
// __block_1559
// __block_1561
_d___pip_5160_1_79___stage___block_26_v_x = _q___pip_5160_1_79___stage___block_26_v_x+_q___pip_5160_1_79___stage___block_26_s_x;

_d___pip_5160_1_79___block_34_tm_x = _q___pip_5160_1_79___block_34_tm_x+_q___pip_5160_1_79___block_40_dt_x;

// __block_1562
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1560
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1563
if (_t___block_1558_y_sel) begin
// __block_1564
// __block_1566
_d___pip_5160_1_79___stage___block_26_v_y = _q___pip_5160_1_79___stage___block_26_v_y+_q___pip_5160_1_79___stage___block_26_s_y;

_d___pip_5160_1_79___block_34_tm_y = _q___pip_5160_1_79___block_34_tm_y+_q___pip_5160_1_79___block_40_dt_y;

// __block_1567
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1565
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1568
if (_t___block_1558_z_sel) begin
// __block_1569
// __block_1571
_d___pip_5160_1_79___stage___block_26_v_z = _q___pip_5160_1_79___stage___block_26_v_z+_q___pip_5160_1_79___stage___block_26_s_z;

_d___pip_5160_1_79___block_34_tm_z = _q___pip_5160_1_79___block_34_tm_z+_q___pip_5160_1_79___block_40_dt_z;

// __block_1572
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1570
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1573
// end of pipeline stage
_d__full_fsm___pip_5160_1_79 = 1;
_d__idx_fsm___pip_5160_1_79 = _t__stall_fsm___pip_5160_1_79 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_79 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 80
(* full_case *)
case (_q__idx_fsm___pip_5160_1_80)
1: begin
// __stage___block_1574
_t___stage___block_1574_tex = (_q___pip_5160_1_80___stage___block_26_v_x)^(_q___pip_5160_1_80___stage___block_26_v_y)^(_q___pip_5160_1_80___stage___block_26_v_z);

_t___stage___block_1574_vnum0 = {_q___pip_5160_1_80___stage___block_26_v_z[0+:2],_q___pip_5160_1_80___stage___block_26_v_y[0+:2],_q___pip_5160_1_80___stage___block_26_v_x[0+:2]};

_t___stage___block_1574_vnum1 = {_q___pip_5160_1_80___stage___block_26_v_z[2+:2],_q___pip_5160_1_80___stage___block_26_v_y[2+:2],_q___pip_5160_1_80___stage___block_26_v_x[2+:2]};

_t___stage___block_1574_vnum2 = {_q___pip_5160_1_80___stage___block_26_v_z[4+:2],_q___pip_5160_1_80___stage___block_26_v_y[4+:2],_q___pip_5160_1_80___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_80___stage___block_6_inside&_w_tile[_t___stage___block_1574_vnum0+:1]&_w_tile[_t___stage___block_1574_vnum1+:1]&_w_tile[_t___stage___block_1574_vnum2+:1]) begin
// __block_1575
// __block_1577
_d___pip_5160_1_80___stage___block_6_clr = _t___stage___block_1574_tex;

_d___pip_5160_1_80___stage___block_6_dist = 136;

_d___pip_5160_1_80___stage___block_6_inside = 1;

// __block_1578
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1576
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1579
_t___block_1579_cmp_yx = _q___pip_5160_1_80___block_34_tm_y-_q___pip_5160_1_80___block_34_tm_x;

_t___block_1579_cmp_zx = _q___pip_5160_1_80___block_34_tm_z-_q___pip_5160_1_80___block_34_tm_x;

_t___block_1579_cmp_zy = _q___pip_5160_1_80___block_34_tm_z-_q___pip_5160_1_80___block_34_tm_y;

_t___block_1579_x_sel = ~_t___block_1579_cmp_yx[20+:1]&&~_t___block_1579_cmp_zx[20+:1];

_t___block_1579_y_sel = _t___block_1579_cmp_yx[20+:1]&&~_t___block_1579_cmp_zy[20+:1];

_t___block_1579_z_sel = _t___block_1579_cmp_zx[20+:1]&&_t___block_1579_cmp_zy[20+:1];

if (_t___block_1579_x_sel) begin
// __block_1580
// __block_1582
_d___pip_5160_1_80___stage___block_26_v_x = _q___pip_5160_1_80___stage___block_26_v_x+_q___pip_5160_1_80___stage___block_26_s_x;

_d___pip_5160_1_80___block_34_tm_x = _q___pip_5160_1_80___block_34_tm_x+_q___pip_5160_1_80___block_40_dt_x;

// __block_1583
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1581
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1584
if (_t___block_1579_y_sel) begin
// __block_1585
// __block_1587
_d___pip_5160_1_80___stage___block_26_v_y = _q___pip_5160_1_80___stage___block_26_v_y+_q___pip_5160_1_80___stage___block_26_s_y;

_d___pip_5160_1_80___block_34_tm_y = _q___pip_5160_1_80___block_34_tm_y+_q___pip_5160_1_80___block_40_dt_y;

// __block_1588
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1586
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1589
if (_t___block_1579_z_sel) begin
// __block_1590
// __block_1592
_d___pip_5160_1_80___stage___block_26_v_z = _q___pip_5160_1_80___stage___block_26_v_z+_q___pip_5160_1_80___stage___block_26_s_z;

_d___pip_5160_1_80___block_34_tm_z = _q___pip_5160_1_80___block_34_tm_z+_q___pip_5160_1_80___block_40_dt_z;

// __block_1593
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1591
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1594
// end of pipeline stage
_d__full_fsm___pip_5160_1_80 = 1;
_d__idx_fsm___pip_5160_1_80 = _t__stall_fsm___pip_5160_1_80 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_80 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 81
(* full_case *)
case (_q__idx_fsm___pip_5160_1_81)
1: begin
// __stage___block_1595
_t___stage___block_1595_tex = (_q___pip_5160_1_81___stage___block_26_v_x)^(_q___pip_5160_1_81___stage___block_26_v_y)^(_q___pip_5160_1_81___stage___block_26_v_z);

_t___stage___block_1595_vnum0 = {_q___pip_5160_1_81___stage___block_26_v_z[0+:2],_q___pip_5160_1_81___stage___block_26_v_y[0+:2],_q___pip_5160_1_81___stage___block_26_v_x[0+:2]};

_t___stage___block_1595_vnum1 = {_q___pip_5160_1_81___stage___block_26_v_z[2+:2],_q___pip_5160_1_81___stage___block_26_v_y[2+:2],_q___pip_5160_1_81___stage___block_26_v_x[2+:2]};

_t___stage___block_1595_vnum2 = {_q___pip_5160_1_81___stage___block_26_v_z[4+:2],_q___pip_5160_1_81___stage___block_26_v_y[4+:2],_q___pip_5160_1_81___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_81___stage___block_6_inside&_w_tile[_t___stage___block_1595_vnum0+:1]&_w_tile[_t___stage___block_1595_vnum1+:1]&_w_tile[_t___stage___block_1595_vnum2+:1]) begin
// __block_1596
// __block_1598
_d___pip_5160_1_81___stage___block_6_clr = _t___stage___block_1595_tex;

_d___pip_5160_1_81___stage___block_6_dist = 138;

_d___pip_5160_1_81___stage___block_6_inside = 1;

// __block_1599
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1597
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1600
_t___block_1600_cmp_yx = _q___pip_5160_1_81___block_34_tm_y-_q___pip_5160_1_81___block_34_tm_x;

_t___block_1600_cmp_zx = _q___pip_5160_1_81___block_34_tm_z-_q___pip_5160_1_81___block_34_tm_x;

_t___block_1600_cmp_zy = _q___pip_5160_1_81___block_34_tm_z-_q___pip_5160_1_81___block_34_tm_y;

_t___block_1600_x_sel = ~_t___block_1600_cmp_yx[20+:1]&&~_t___block_1600_cmp_zx[20+:1];

_t___block_1600_y_sel = _t___block_1600_cmp_yx[20+:1]&&~_t___block_1600_cmp_zy[20+:1];

_t___block_1600_z_sel = _t___block_1600_cmp_zx[20+:1]&&_t___block_1600_cmp_zy[20+:1];

if (_t___block_1600_x_sel) begin
// __block_1601
// __block_1603
_d___pip_5160_1_81___stage___block_26_v_x = _q___pip_5160_1_81___stage___block_26_v_x+_q___pip_5160_1_81___stage___block_26_s_x;

_d___pip_5160_1_81___block_34_tm_x = _q___pip_5160_1_81___block_34_tm_x+_q___pip_5160_1_81___block_40_dt_x;

// __block_1604
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1602
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1605
if (_t___block_1600_y_sel) begin
// __block_1606
// __block_1608
_d___pip_5160_1_81___stage___block_26_v_y = _q___pip_5160_1_81___stage___block_26_v_y+_q___pip_5160_1_81___stage___block_26_s_y;

_d___pip_5160_1_81___block_34_tm_y = _q___pip_5160_1_81___block_34_tm_y+_q___pip_5160_1_81___block_40_dt_y;

// __block_1609
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1607
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1610
if (_t___block_1600_z_sel) begin
// __block_1611
// __block_1613
_d___pip_5160_1_81___stage___block_26_v_z = _q___pip_5160_1_81___stage___block_26_v_z+_q___pip_5160_1_81___stage___block_26_s_z;

_d___pip_5160_1_81___block_34_tm_z = _q___pip_5160_1_81___block_34_tm_z+_q___pip_5160_1_81___block_40_dt_z;

// __block_1614
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1612
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1615
// end of pipeline stage
_d__full_fsm___pip_5160_1_81 = 1;
_d__idx_fsm___pip_5160_1_81 = _t__stall_fsm___pip_5160_1_81 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_81 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 82
(* full_case *)
case (_q__idx_fsm___pip_5160_1_82)
1: begin
// __stage___block_1616
_t___stage___block_1616_tex = (_q___pip_5160_1_82___stage___block_26_v_x)^(_q___pip_5160_1_82___stage___block_26_v_y)^(_q___pip_5160_1_82___stage___block_26_v_z);

_t___stage___block_1616_vnum0 = {_q___pip_5160_1_82___stage___block_26_v_z[0+:2],_q___pip_5160_1_82___stage___block_26_v_y[0+:2],_q___pip_5160_1_82___stage___block_26_v_x[0+:2]};

_t___stage___block_1616_vnum1 = {_q___pip_5160_1_82___stage___block_26_v_z[2+:2],_q___pip_5160_1_82___stage___block_26_v_y[2+:2],_q___pip_5160_1_82___stage___block_26_v_x[2+:2]};

_t___stage___block_1616_vnum2 = {_q___pip_5160_1_82___stage___block_26_v_z[4+:2],_q___pip_5160_1_82___stage___block_26_v_y[4+:2],_q___pip_5160_1_82___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_82___stage___block_6_inside&_w_tile[_t___stage___block_1616_vnum0+:1]&_w_tile[_t___stage___block_1616_vnum1+:1]&_w_tile[_t___stage___block_1616_vnum2+:1]) begin
// __block_1617
// __block_1619
_d___pip_5160_1_82___stage___block_6_clr = _t___stage___block_1616_tex;

_d___pip_5160_1_82___stage___block_6_dist = 140;

_d___pip_5160_1_82___stage___block_6_inside = 1;

// __block_1620
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1618
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1621
_t___block_1621_cmp_yx = _q___pip_5160_1_82___block_34_tm_y-_q___pip_5160_1_82___block_34_tm_x;

_t___block_1621_cmp_zx = _q___pip_5160_1_82___block_34_tm_z-_q___pip_5160_1_82___block_34_tm_x;

_t___block_1621_cmp_zy = _q___pip_5160_1_82___block_34_tm_z-_q___pip_5160_1_82___block_34_tm_y;

_t___block_1621_x_sel = ~_t___block_1621_cmp_yx[20+:1]&&~_t___block_1621_cmp_zx[20+:1];

_t___block_1621_y_sel = _t___block_1621_cmp_yx[20+:1]&&~_t___block_1621_cmp_zy[20+:1];

_t___block_1621_z_sel = _t___block_1621_cmp_zx[20+:1]&&_t___block_1621_cmp_zy[20+:1];

if (_t___block_1621_x_sel) begin
// __block_1622
// __block_1624
_d___pip_5160_1_82___stage___block_26_v_x = _q___pip_5160_1_82___stage___block_26_v_x+_q___pip_5160_1_82___stage___block_26_s_x;

_d___pip_5160_1_82___block_34_tm_x = _q___pip_5160_1_82___block_34_tm_x+_q___pip_5160_1_82___block_40_dt_x;

// __block_1625
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1623
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1626
if (_t___block_1621_y_sel) begin
// __block_1627
// __block_1629
_d___pip_5160_1_82___stage___block_26_v_y = _q___pip_5160_1_82___stage___block_26_v_y+_q___pip_5160_1_82___stage___block_26_s_y;

_d___pip_5160_1_82___block_34_tm_y = _q___pip_5160_1_82___block_34_tm_y+_q___pip_5160_1_82___block_40_dt_y;

// __block_1630
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1628
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1631
if (_t___block_1621_z_sel) begin
// __block_1632
// __block_1634
_d___pip_5160_1_82___stage___block_26_v_z = _q___pip_5160_1_82___stage___block_26_v_z+_q___pip_5160_1_82___stage___block_26_s_z;

_d___pip_5160_1_82___block_34_tm_z = _q___pip_5160_1_82___block_34_tm_z+_q___pip_5160_1_82___block_40_dt_z;

// __block_1635
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1633
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1636
// end of pipeline stage
_d__full_fsm___pip_5160_1_82 = 1;
_d__idx_fsm___pip_5160_1_82 = _t__stall_fsm___pip_5160_1_82 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_82 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 83
(* full_case *)
case (_q__idx_fsm___pip_5160_1_83)
1: begin
// __stage___block_1637
_t___stage___block_1637_tex = (_q___pip_5160_1_83___stage___block_26_v_x)^(_q___pip_5160_1_83___stage___block_26_v_y)^(_q___pip_5160_1_83___stage___block_26_v_z);

_t___stage___block_1637_vnum0 = {_q___pip_5160_1_83___stage___block_26_v_z[0+:2],_q___pip_5160_1_83___stage___block_26_v_y[0+:2],_q___pip_5160_1_83___stage___block_26_v_x[0+:2]};

_t___stage___block_1637_vnum1 = {_q___pip_5160_1_83___stage___block_26_v_z[2+:2],_q___pip_5160_1_83___stage___block_26_v_y[2+:2],_q___pip_5160_1_83___stage___block_26_v_x[2+:2]};

_t___stage___block_1637_vnum2 = {_q___pip_5160_1_83___stage___block_26_v_z[4+:2],_q___pip_5160_1_83___stage___block_26_v_y[4+:2],_q___pip_5160_1_83___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_83___stage___block_6_inside&_w_tile[_t___stage___block_1637_vnum0+:1]&_w_tile[_t___stage___block_1637_vnum1+:1]&_w_tile[_t___stage___block_1637_vnum2+:1]) begin
// __block_1638
// __block_1640
_d___pip_5160_1_83___stage___block_6_clr = _t___stage___block_1637_tex;

_d___pip_5160_1_83___stage___block_6_dist = 141;

_d___pip_5160_1_83___stage___block_6_inside = 1;

// __block_1641
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1639
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1642
_t___block_1642_cmp_yx = _q___pip_5160_1_83___block_34_tm_y-_q___pip_5160_1_83___block_34_tm_x;

_t___block_1642_cmp_zx = _q___pip_5160_1_83___block_34_tm_z-_q___pip_5160_1_83___block_34_tm_x;

_t___block_1642_cmp_zy = _q___pip_5160_1_83___block_34_tm_z-_q___pip_5160_1_83___block_34_tm_y;

_t___block_1642_x_sel = ~_t___block_1642_cmp_yx[20+:1]&&~_t___block_1642_cmp_zx[20+:1];

_t___block_1642_y_sel = _t___block_1642_cmp_yx[20+:1]&&~_t___block_1642_cmp_zy[20+:1];

_t___block_1642_z_sel = _t___block_1642_cmp_zx[20+:1]&&_t___block_1642_cmp_zy[20+:1];

if (_t___block_1642_x_sel) begin
// __block_1643
// __block_1645
_d___pip_5160_1_83___stage___block_26_v_x = _q___pip_5160_1_83___stage___block_26_v_x+_q___pip_5160_1_83___stage___block_26_s_x;

_d___pip_5160_1_83___block_34_tm_x = _q___pip_5160_1_83___block_34_tm_x+_q___pip_5160_1_83___block_40_dt_x;

// __block_1646
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1644
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1647
if (_t___block_1642_y_sel) begin
// __block_1648
// __block_1650
_d___pip_5160_1_83___stage___block_26_v_y = _q___pip_5160_1_83___stage___block_26_v_y+_q___pip_5160_1_83___stage___block_26_s_y;

_d___pip_5160_1_83___block_34_tm_y = _q___pip_5160_1_83___block_34_tm_y+_q___pip_5160_1_83___block_40_dt_y;

// __block_1651
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1649
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1652
if (_t___block_1642_z_sel) begin
// __block_1653
// __block_1655
_d___pip_5160_1_83___stage___block_26_v_z = _q___pip_5160_1_83___stage___block_26_v_z+_q___pip_5160_1_83___stage___block_26_s_z;

_d___pip_5160_1_83___block_34_tm_z = _q___pip_5160_1_83___block_34_tm_z+_q___pip_5160_1_83___block_40_dt_z;

// __block_1656
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1654
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1657
// end of pipeline stage
_d__full_fsm___pip_5160_1_83 = 1;
_d__idx_fsm___pip_5160_1_83 = _t__stall_fsm___pip_5160_1_83 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_83 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 84
(* full_case *)
case (_q__idx_fsm___pip_5160_1_84)
1: begin
// __stage___block_1658
_t___stage___block_1658_tex = (_q___pip_5160_1_84___stage___block_26_v_x)^(_q___pip_5160_1_84___stage___block_26_v_y)^(_q___pip_5160_1_84___stage___block_26_v_z);

_t___stage___block_1658_vnum0 = {_q___pip_5160_1_84___stage___block_26_v_z[0+:2],_q___pip_5160_1_84___stage___block_26_v_y[0+:2],_q___pip_5160_1_84___stage___block_26_v_x[0+:2]};

_t___stage___block_1658_vnum1 = {_q___pip_5160_1_84___stage___block_26_v_z[2+:2],_q___pip_5160_1_84___stage___block_26_v_y[2+:2],_q___pip_5160_1_84___stage___block_26_v_x[2+:2]};

_t___stage___block_1658_vnum2 = {_q___pip_5160_1_84___stage___block_26_v_z[4+:2],_q___pip_5160_1_84___stage___block_26_v_y[4+:2],_q___pip_5160_1_84___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_84___stage___block_6_inside&_w_tile[_t___stage___block_1658_vnum0+:1]&_w_tile[_t___stage___block_1658_vnum1+:1]&_w_tile[_t___stage___block_1658_vnum2+:1]) begin
// __block_1659
// __block_1661
_d___pip_5160_1_84___stage___block_6_clr = _t___stage___block_1658_tex;

_d___pip_5160_1_84___stage___block_6_dist = 143;

_d___pip_5160_1_84___stage___block_6_inside = 1;

// __block_1662
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1660
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1663
_t___block_1663_cmp_yx = _q___pip_5160_1_84___block_34_tm_y-_q___pip_5160_1_84___block_34_tm_x;

_t___block_1663_cmp_zx = _q___pip_5160_1_84___block_34_tm_z-_q___pip_5160_1_84___block_34_tm_x;

_t___block_1663_cmp_zy = _q___pip_5160_1_84___block_34_tm_z-_q___pip_5160_1_84___block_34_tm_y;

_t___block_1663_x_sel = ~_t___block_1663_cmp_yx[20+:1]&&~_t___block_1663_cmp_zx[20+:1];

_t___block_1663_y_sel = _t___block_1663_cmp_yx[20+:1]&&~_t___block_1663_cmp_zy[20+:1];

_t___block_1663_z_sel = _t___block_1663_cmp_zx[20+:1]&&_t___block_1663_cmp_zy[20+:1];

if (_t___block_1663_x_sel) begin
// __block_1664
// __block_1666
_d___pip_5160_1_84___stage___block_26_v_x = _q___pip_5160_1_84___stage___block_26_v_x+_q___pip_5160_1_84___stage___block_26_s_x;

_d___pip_5160_1_84___block_34_tm_x = _q___pip_5160_1_84___block_34_tm_x+_q___pip_5160_1_84___block_40_dt_x;

// __block_1667
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1665
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1668
if (_t___block_1663_y_sel) begin
// __block_1669
// __block_1671
_d___pip_5160_1_84___stage___block_26_v_y = _q___pip_5160_1_84___stage___block_26_v_y+_q___pip_5160_1_84___stage___block_26_s_y;

_d___pip_5160_1_84___block_34_tm_y = _q___pip_5160_1_84___block_34_tm_y+_q___pip_5160_1_84___block_40_dt_y;

// __block_1672
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1670
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1673
if (_t___block_1663_z_sel) begin
// __block_1674
// __block_1676
_d___pip_5160_1_84___stage___block_26_v_z = _q___pip_5160_1_84___stage___block_26_v_z+_q___pip_5160_1_84___stage___block_26_s_z;

_d___pip_5160_1_84___block_34_tm_z = _q___pip_5160_1_84___block_34_tm_z+_q___pip_5160_1_84___block_40_dt_z;

// __block_1677
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1675
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1678
// end of pipeline stage
_d__full_fsm___pip_5160_1_84 = 1;
_d__idx_fsm___pip_5160_1_84 = _t__stall_fsm___pip_5160_1_84 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_84 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 85
(* full_case *)
case (_q__idx_fsm___pip_5160_1_85)
1: begin
// __stage___block_1679
_t___stage___block_1679_tex = (_q___pip_5160_1_85___stage___block_26_v_x)^(_q___pip_5160_1_85___stage___block_26_v_y)^(_q___pip_5160_1_85___stage___block_26_v_z);

_t___stage___block_1679_vnum0 = {_q___pip_5160_1_85___stage___block_26_v_z[0+:2],_q___pip_5160_1_85___stage___block_26_v_y[0+:2],_q___pip_5160_1_85___stage___block_26_v_x[0+:2]};

_t___stage___block_1679_vnum1 = {_q___pip_5160_1_85___stage___block_26_v_z[2+:2],_q___pip_5160_1_85___stage___block_26_v_y[2+:2],_q___pip_5160_1_85___stage___block_26_v_x[2+:2]};

_t___stage___block_1679_vnum2 = {_q___pip_5160_1_85___stage___block_26_v_z[4+:2],_q___pip_5160_1_85___stage___block_26_v_y[4+:2],_q___pip_5160_1_85___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_85___stage___block_6_inside&_w_tile[_t___stage___block_1679_vnum0+:1]&_w_tile[_t___stage___block_1679_vnum1+:1]&_w_tile[_t___stage___block_1679_vnum2+:1]) begin
// __block_1680
// __block_1682
_d___pip_5160_1_85___stage___block_6_clr = _t___stage___block_1679_tex;

_d___pip_5160_1_85___stage___block_6_dist = 145;

_d___pip_5160_1_85___stage___block_6_inside = 1;

// __block_1683
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1681
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1684
_t___block_1684_cmp_yx = _q___pip_5160_1_85___block_34_tm_y-_q___pip_5160_1_85___block_34_tm_x;

_t___block_1684_cmp_zx = _q___pip_5160_1_85___block_34_tm_z-_q___pip_5160_1_85___block_34_tm_x;

_t___block_1684_cmp_zy = _q___pip_5160_1_85___block_34_tm_z-_q___pip_5160_1_85___block_34_tm_y;

_t___block_1684_x_sel = ~_t___block_1684_cmp_yx[20+:1]&&~_t___block_1684_cmp_zx[20+:1];

_t___block_1684_y_sel = _t___block_1684_cmp_yx[20+:1]&&~_t___block_1684_cmp_zy[20+:1];

_t___block_1684_z_sel = _t___block_1684_cmp_zx[20+:1]&&_t___block_1684_cmp_zy[20+:1];

if (_t___block_1684_x_sel) begin
// __block_1685
// __block_1687
_d___pip_5160_1_85___stage___block_26_v_x = _q___pip_5160_1_85___stage___block_26_v_x+_q___pip_5160_1_85___stage___block_26_s_x;

_d___pip_5160_1_85___block_34_tm_x = _q___pip_5160_1_85___block_34_tm_x+_q___pip_5160_1_85___block_40_dt_x;

// __block_1688
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1686
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1689
if (_t___block_1684_y_sel) begin
// __block_1690
// __block_1692
_d___pip_5160_1_85___stage___block_26_v_y = _q___pip_5160_1_85___stage___block_26_v_y+_q___pip_5160_1_85___stage___block_26_s_y;

_d___pip_5160_1_85___block_34_tm_y = _q___pip_5160_1_85___block_34_tm_y+_q___pip_5160_1_85___block_40_dt_y;

// __block_1693
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1691
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1694
if (_t___block_1684_z_sel) begin
// __block_1695
// __block_1697
_d___pip_5160_1_85___stage___block_26_v_z = _q___pip_5160_1_85___stage___block_26_v_z+_q___pip_5160_1_85___stage___block_26_s_z;

_d___pip_5160_1_85___block_34_tm_z = _q___pip_5160_1_85___block_34_tm_z+_q___pip_5160_1_85___block_40_dt_z;

// __block_1698
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1696
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1699
// end of pipeline stage
_d__full_fsm___pip_5160_1_85 = 1;
_d__idx_fsm___pip_5160_1_85 = _t__stall_fsm___pip_5160_1_85 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_85 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 86
(* full_case *)
case (_q__idx_fsm___pip_5160_1_86)
1: begin
// __stage___block_1700
_t___stage___block_1700_tex = (_q___pip_5160_1_86___stage___block_26_v_x)^(_q___pip_5160_1_86___stage___block_26_v_y)^(_q___pip_5160_1_86___stage___block_26_v_z);

_t___stage___block_1700_vnum0 = {_q___pip_5160_1_86___stage___block_26_v_z[0+:2],_q___pip_5160_1_86___stage___block_26_v_y[0+:2],_q___pip_5160_1_86___stage___block_26_v_x[0+:2]};

_t___stage___block_1700_vnum1 = {_q___pip_5160_1_86___stage___block_26_v_z[2+:2],_q___pip_5160_1_86___stage___block_26_v_y[2+:2],_q___pip_5160_1_86___stage___block_26_v_x[2+:2]};

_t___stage___block_1700_vnum2 = {_q___pip_5160_1_86___stage___block_26_v_z[4+:2],_q___pip_5160_1_86___stage___block_26_v_y[4+:2],_q___pip_5160_1_86___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_86___stage___block_6_inside&_w_tile[_t___stage___block_1700_vnum0+:1]&_w_tile[_t___stage___block_1700_vnum1+:1]&_w_tile[_t___stage___block_1700_vnum2+:1]) begin
// __block_1701
// __block_1703
_d___pip_5160_1_86___stage___block_6_clr = _t___stage___block_1700_tex;

_d___pip_5160_1_86___stage___block_6_dist = 147;

_d___pip_5160_1_86___stage___block_6_inside = 1;

// __block_1704
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1702
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1705
_t___block_1705_cmp_yx = _q___pip_5160_1_86___block_34_tm_y-_q___pip_5160_1_86___block_34_tm_x;

_t___block_1705_cmp_zx = _q___pip_5160_1_86___block_34_tm_z-_q___pip_5160_1_86___block_34_tm_x;

_t___block_1705_cmp_zy = _q___pip_5160_1_86___block_34_tm_z-_q___pip_5160_1_86___block_34_tm_y;

_t___block_1705_x_sel = ~_t___block_1705_cmp_yx[20+:1]&&~_t___block_1705_cmp_zx[20+:1];

_t___block_1705_y_sel = _t___block_1705_cmp_yx[20+:1]&&~_t___block_1705_cmp_zy[20+:1];

_t___block_1705_z_sel = _t___block_1705_cmp_zx[20+:1]&&_t___block_1705_cmp_zy[20+:1];

if (_t___block_1705_x_sel) begin
// __block_1706
// __block_1708
_d___pip_5160_1_86___stage___block_26_v_x = _q___pip_5160_1_86___stage___block_26_v_x+_q___pip_5160_1_86___stage___block_26_s_x;

_d___pip_5160_1_86___block_34_tm_x = _q___pip_5160_1_86___block_34_tm_x+_q___pip_5160_1_86___block_40_dt_x;

// __block_1709
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1707
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1710
if (_t___block_1705_y_sel) begin
// __block_1711
// __block_1713
_d___pip_5160_1_86___stage___block_26_v_y = _q___pip_5160_1_86___stage___block_26_v_y+_q___pip_5160_1_86___stage___block_26_s_y;

_d___pip_5160_1_86___block_34_tm_y = _q___pip_5160_1_86___block_34_tm_y+_q___pip_5160_1_86___block_40_dt_y;

// __block_1714
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1712
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1715
if (_t___block_1705_z_sel) begin
// __block_1716
// __block_1718
_d___pip_5160_1_86___stage___block_26_v_z = _q___pip_5160_1_86___stage___block_26_v_z+_q___pip_5160_1_86___stage___block_26_s_z;

_d___pip_5160_1_86___block_34_tm_z = _q___pip_5160_1_86___block_34_tm_z+_q___pip_5160_1_86___block_40_dt_z;

// __block_1719
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1717
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1720
// end of pipeline stage
_d__full_fsm___pip_5160_1_86 = 1;
_d__idx_fsm___pip_5160_1_86 = _t__stall_fsm___pip_5160_1_86 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_86 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 87
(* full_case *)
case (_q__idx_fsm___pip_5160_1_87)
1: begin
// __stage___block_1721
_t___stage___block_1721_tex = (_q___pip_5160_1_87___stage___block_26_v_x)^(_q___pip_5160_1_87___stage___block_26_v_y)^(_q___pip_5160_1_87___stage___block_26_v_z);

_t___stage___block_1721_vnum0 = {_q___pip_5160_1_87___stage___block_26_v_z[0+:2],_q___pip_5160_1_87___stage___block_26_v_y[0+:2],_q___pip_5160_1_87___stage___block_26_v_x[0+:2]};

_t___stage___block_1721_vnum1 = {_q___pip_5160_1_87___stage___block_26_v_z[2+:2],_q___pip_5160_1_87___stage___block_26_v_y[2+:2],_q___pip_5160_1_87___stage___block_26_v_x[2+:2]};

_t___stage___block_1721_vnum2 = {_q___pip_5160_1_87___stage___block_26_v_z[4+:2],_q___pip_5160_1_87___stage___block_26_v_y[4+:2],_q___pip_5160_1_87___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_87___stage___block_6_inside&_w_tile[_t___stage___block_1721_vnum0+:1]&_w_tile[_t___stage___block_1721_vnum1+:1]&_w_tile[_t___stage___block_1721_vnum2+:1]) begin
// __block_1722
// __block_1724
_d___pip_5160_1_87___stage___block_6_clr = _t___stage___block_1721_tex;

_d___pip_5160_1_87___stage___block_6_dist = 149;

_d___pip_5160_1_87___stage___block_6_inside = 1;

// __block_1725
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1723
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1726
_t___block_1726_cmp_yx = _q___pip_5160_1_87___block_34_tm_y-_q___pip_5160_1_87___block_34_tm_x;

_t___block_1726_cmp_zx = _q___pip_5160_1_87___block_34_tm_z-_q___pip_5160_1_87___block_34_tm_x;

_t___block_1726_cmp_zy = _q___pip_5160_1_87___block_34_tm_z-_q___pip_5160_1_87___block_34_tm_y;

_t___block_1726_x_sel = ~_t___block_1726_cmp_yx[20+:1]&&~_t___block_1726_cmp_zx[20+:1];

_t___block_1726_y_sel = _t___block_1726_cmp_yx[20+:1]&&~_t___block_1726_cmp_zy[20+:1];

_t___block_1726_z_sel = _t___block_1726_cmp_zx[20+:1]&&_t___block_1726_cmp_zy[20+:1];

if (_t___block_1726_x_sel) begin
// __block_1727
// __block_1729
_d___pip_5160_1_87___stage___block_26_v_x = _q___pip_5160_1_87___stage___block_26_v_x+_q___pip_5160_1_87___stage___block_26_s_x;

_d___pip_5160_1_87___block_34_tm_x = _q___pip_5160_1_87___block_34_tm_x+_q___pip_5160_1_87___block_40_dt_x;

// __block_1730
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1728
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1731
if (_t___block_1726_y_sel) begin
// __block_1732
// __block_1734
_d___pip_5160_1_87___stage___block_26_v_y = _q___pip_5160_1_87___stage___block_26_v_y+_q___pip_5160_1_87___stage___block_26_s_y;

_d___pip_5160_1_87___block_34_tm_y = _q___pip_5160_1_87___block_34_tm_y+_q___pip_5160_1_87___block_40_dt_y;

// __block_1735
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1733
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1736
if (_t___block_1726_z_sel) begin
// __block_1737
// __block_1739
_d___pip_5160_1_87___stage___block_26_v_z = _q___pip_5160_1_87___stage___block_26_v_z+_q___pip_5160_1_87___stage___block_26_s_z;

_d___pip_5160_1_87___block_34_tm_z = _q___pip_5160_1_87___block_34_tm_z+_q___pip_5160_1_87___block_40_dt_z;

// __block_1740
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1738
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1741
// end of pipeline stage
_d__full_fsm___pip_5160_1_87 = 1;
_d__idx_fsm___pip_5160_1_87 = _t__stall_fsm___pip_5160_1_87 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_87 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 88
(* full_case *)
case (_q__idx_fsm___pip_5160_1_88)
1: begin
// __stage___block_1742
_t___stage___block_1742_tex = (_q___pip_5160_1_88___stage___block_26_v_x)^(_q___pip_5160_1_88___stage___block_26_v_y)^(_q___pip_5160_1_88___stage___block_26_v_z);

_t___stage___block_1742_vnum0 = {_q___pip_5160_1_88___stage___block_26_v_z[0+:2],_q___pip_5160_1_88___stage___block_26_v_y[0+:2],_q___pip_5160_1_88___stage___block_26_v_x[0+:2]};

_t___stage___block_1742_vnum1 = {_q___pip_5160_1_88___stage___block_26_v_z[2+:2],_q___pip_5160_1_88___stage___block_26_v_y[2+:2],_q___pip_5160_1_88___stage___block_26_v_x[2+:2]};

_t___stage___block_1742_vnum2 = {_q___pip_5160_1_88___stage___block_26_v_z[4+:2],_q___pip_5160_1_88___stage___block_26_v_y[4+:2],_q___pip_5160_1_88___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_88___stage___block_6_inside&_w_tile[_t___stage___block_1742_vnum0+:1]&_w_tile[_t___stage___block_1742_vnum1+:1]&_w_tile[_t___stage___block_1742_vnum2+:1]) begin
// __block_1743
// __block_1745
_d___pip_5160_1_88___stage___block_6_clr = _t___stage___block_1742_tex;

_d___pip_5160_1_88___stage___block_6_dist = 151;

_d___pip_5160_1_88___stage___block_6_inside = 1;

// __block_1746
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1744
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1747
_t___block_1747_cmp_yx = _q___pip_5160_1_88___block_34_tm_y-_q___pip_5160_1_88___block_34_tm_x;

_t___block_1747_cmp_zx = _q___pip_5160_1_88___block_34_tm_z-_q___pip_5160_1_88___block_34_tm_x;

_t___block_1747_cmp_zy = _q___pip_5160_1_88___block_34_tm_z-_q___pip_5160_1_88___block_34_tm_y;

_t___block_1747_x_sel = ~_t___block_1747_cmp_yx[20+:1]&&~_t___block_1747_cmp_zx[20+:1];

_t___block_1747_y_sel = _t___block_1747_cmp_yx[20+:1]&&~_t___block_1747_cmp_zy[20+:1];

_t___block_1747_z_sel = _t___block_1747_cmp_zx[20+:1]&&_t___block_1747_cmp_zy[20+:1];

if (_t___block_1747_x_sel) begin
// __block_1748
// __block_1750
_d___pip_5160_1_88___stage___block_26_v_x = _q___pip_5160_1_88___stage___block_26_v_x+_q___pip_5160_1_88___stage___block_26_s_x;

_d___pip_5160_1_88___block_34_tm_x = _q___pip_5160_1_88___block_34_tm_x+_q___pip_5160_1_88___block_40_dt_x;

// __block_1751
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1749
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1752
if (_t___block_1747_y_sel) begin
// __block_1753
// __block_1755
_d___pip_5160_1_88___stage___block_26_v_y = _q___pip_5160_1_88___stage___block_26_v_y+_q___pip_5160_1_88___stage___block_26_s_y;

_d___pip_5160_1_88___block_34_tm_y = _q___pip_5160_1_88___block_34_tm_y+_q___pip_5160_1_88___block_40_dt_y;

// __block_1756
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1754
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1757
if (_t___block_1747_z_sel) begin
// __block_1758
// __block_1760
_d___pip_5160_1_88___stage___block_26_v_z = _q___pip_5160_1_88___stage___block_26_v_z+_q___pip_5160_1_88___stage___block_26_s_z;

_d___pip_5160_1_88___block_34_tm_z = _q___pip_5160_1_88___block_34_tm_z+_q___pip_5160_1_88___block_40_dt_z;

// __block_1761
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1759
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1762
// end of pipeline stage
_d__full_fsm___pip_5160_1_88 = 1;
_d__idx_fsm___pip_5160_1_88 = _t__stall_fsm___pip_5160_1_88 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_88 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 89
(* full_case *)
case (_q__idx_fsm___pip_5160_1_89)
1: begin
// __stage___block_1763
_t___stage___block_1763_tex = (_q___pip_5160_1_89___stage___block_26_v_x)^(_q___pip_5160_1_89___stage___block_26_v_y)^(_q___pip_5160_1_89___stage___block_26_v_z);

_t___stage___block_1763_vnum0 = {_q___pip_5160_1_89___stage___block_26_v_z[0+:2],_q___pip_5160_1_89___stage___block_26_v_y[0+:2],_q___pip_5160_1_89___stage___block_26_v_x[0+:2]};

_t___stage___block_1763_vnum1 = {_q___pip_5160_1_89___stage___block_26_v_z[2+:2],_q___pip_5160_1_89___stage___block_26_v_y[2+:2],_q___pip_5160_1_89___stage___block_26_v_x[2+:2]};

_t___stage___block_1763_vnum2 = {_q___pip_5160_1_89___stage___block_26_v_z[4+:2],_q___pip_5160_1_89___stage___block_26_v_y[4+:2],_q___pip_5160_1_89___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_89___stage___block_6_inside&_w_tile[_t___stage___block_1763_vnum0+:1]&_w_tile[_t___stage___block_1763_vnum1+:1]&_w_tile[_t___stage___block_1763_vnum2+:1]) begin
// __block_1764
// __block_1766
_d___pip_5160_1_89___stage___block_6_clr = _t___stage___block_1763_tex;

_d___pip_5160_1_89___stage___block_6_dist = 153;

_d___pip_5160_1_89___stage___block_6_inside = 1;

// __block_1767
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1765
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1768
_t___block_1768_cmp_yx = _q___pip_5160_1_89___block_34_tm_y-_q___pip_5160_1_89___block_34_tm_x;

_t___block_1768_cmp_zx = _q___pip_5160_1_89___block_34_tm_z-_q___pip_5160_1_89___block_34_tm_x;

_t___block_1768_cmp_zy = _q___pip_5160_1_89___block_34_tm_z-_q___pip_5160_1_89___block_34_tm_y;

_t___block_1768_x_sel = ~_t___block_1768_cmp_yx[20+:1]&&~_t___block_1768_cmp_zx[20+:1];

_t___block_1768_y_sel = _t___block_1768_cmp_yx[20+:1]&&~_t___block_1768_cmp_zy[20+:1];

_t___block_1768_z_sel = _t___block_1768_cmp_zx[20+:1]&&_t___block_1768_cmp_zy[20+:1];

if (_t___block_1768_x_sel) begin
// __block_1769
// __block_1771
_d___pip_5160_1_89___stage___block_26_v_x = _q___pip_5160_1_89___stage___block_26_v_x+_q___pip_5160_1_89___stage___block_26_s_x;

_d___pip_5160_1_89___block_34_tm_x = _q___pip_5160_1_89___block_34_tm_x+_q___pip_5160_1_89___block_40_dt_x;

// __block_1772
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1770
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1773
if (_t___block_1768_y_sel) begin
// __block_1774
// __block_1776
_d___pip_5160_1_89___stage___block_26_v_y = _q___pip_5160_1_89___stage___block_26_v_y+_q___pip_5160_1_89___stage___block_26_s_y;

_d___pip_5160_1_89___block_34_tm_y = _q___pip_5160_1_89___block_34_tm_y+_q___pip_5160_1_89___block_40_dt_y;

// __block_1777
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1775
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1778
if (_t___block_1768_z_sel) begin
// __block_1779
// __block_1781
_d___pip_5160_1_89___stage___block_26_v_z = _q___pip_5160_1_89___stage___block_26_v_z+_q___pip_5160_1_89___stage___block_26_s_z;

_d___pip_5160_1_89___block_34_tm_z = _q___pip_5160_1_89___block_34_tm_z+_q___pip_5160_1_89___block_40_dt_z;

// __block_1782
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1780
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1783
// end of pipeline stage
_d__full_fsm___pip_5160_1_89 = 1;
_d__idx_fsm___pip_5160_1_89 = _t__stall_fsm___pip_5160_1_89 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_89 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 90
(* full_case *)
case (_q__idx_fsm___pip_5160_1_90)
1: begin
// __stage___block_1784
_t___stage___block_1784_tex = (_q___pip_5160_1_90___stage___block_26_v_x)^(_q___pip_5160_1_90___stage___block_26_v_y)^(_q___pip_5160_1_90___stage___block_26_v_z);

_t___stage___block_1784_vnum0 = {_q___pip_5160_1_90___stage___block_26_v_z[0+:2],_q___pip_5160_1_90___stage___block_26_v_y[0+:2],_q___pip_5160_1_90___stage___block_26_v_x[0+:2]};

_t___stage___block_1784_vnum1 = {_q___pip_5160_1_90___stage___block_26_v_z[2+:2],_q___pip_5160_1_90___stage___block_26_v_y[2+:2],_q___pip_5160_1_90___stage___block_26_v_x[2+:2]};

_t___stage___block_1784_vnum2 = {_q___pip_5160_1_90___stage___block_26_v_z[4+:2],_q___pip_5160_1_90___stage___block_26_v_y[4+:2],_q___pip_5160_1_90___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_90___stage___block_6_inside&_w_tile[_t___stage___block_1784_vnum0+:1]&_w_tile[_t___stage___block_1784_vnum1+:1]&_w_tile[_t___stage___block_1784_vnum2+:1]) begin
// __block_1785
// __block_1787
_d___pip_5160_1_90___stage___block_6_clr = _t___stage___block_1784_tex;

_d___pip_5160_1_90___stage___block_6_dist = 154;

_d___pip_5160_1_90___stage___block_6_inside = 1;

// __block_1788
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1786
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1789
_t___block_1789_cmp_yx = _q___pip_5160_1_90___block_34_tm_y-_q___pip_5160_1_90___block_34_tm_x;

_t___block_1789_cmp_zx = _q___pip_5160_1_90___block_34_tm_z-_q___pip_5160_1_90___block_34_tm_x;

_t___block_1789_cmp_zy = _q___pip_5160_1_90___block_34_tm_z-_q___pip_5160_1_90___block_34_tm_y;

_t___block_1789_x_sel = ~_t___block_1789_cmp_yx[20+:1]&&~_t___block_1789_cmp_zx[20+:1];

_t___block_1789_y_sel = _t___block_1789_cmp_yx[20+:1]&&~_t___block_1789_cmp_zy[20+:1];

_t___block_1789_z_sel = _t___block_1789_cmp_zx[20+:1]&&_t___block_1789_cmp_zy[20+:1];

if (_t___block_1789_x_sel) begin
// __block_1790
// __block_1792
_d___pip_5160_1_90___stage___block_26_v_x = _q___pip_5160_1_90___stage___block_26_v_x+_q___pip_5160_1_90___stage___block_26_s_x;

_d___pip_5160_1_90___block_34_tm_x = _q___pip_5160_1_90___block_34_tm_x+_q___pip_5160_1_90___block_40_dt_x;

// __block_1793
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1791
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1794
if (_t___block_1789_y_sel) begin
// __block_1795
// __block_1797
_d___pip_5160_1_90___stage___block_26_v_y = _q___pip_5160_1_90___stage___block_26_v_y+_q___pip_5160_1_90___stage___block_26_s_y;

_d___pip_5160_1_90___block_34_tm_y = _q___pip_5160_1_90___block_34_tm_y+_q___pip_5160_1_90___block_40_dt_y;

// __block_1798
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1796
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1799
if (_t___block_1789_z_sel) begin
// __block_1800
// __block_1802
_d___pip_5160_1_90___stage___block_26_v_z = _q___pip_5160_1_90___stage___block_26_v_z+_q___pip_5160_1_90___stage___block_26_s_z;

_d___pip_5160_1_90___block_34_tm_z = _q___pip_5160_1_90___block_34_tm_z+_q___pip_5160_1_90___block_40_dt_z;

// __block_1803
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1801
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1804
// end of pipeline stage
_d__full_fsm___pip_5160_1_90 = 1;
_d__idx_fsm___pip_5160_1_90 = _t__stall_fsm___pip_5160_1_90 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_90 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 91
(* full_case *)
case (_q__idx_fsm___pip_5160_1_91)
1: begin
// __stage___block_1805
_t___stage___block_1805_tex = (_q___pip_5160_1_91___stage___block_26_v_x)^(_q___pip_5160_1_91___stage___block_26_v_y)^(_q___pip_5160_1_91___stage___block_26_v_z);

_t___stage___block_1805_vnum0 = {_q___pip_5160_1_91___stage___block_26_v_z[0+:2],_q___pip_5160_1_91___stage___block_26_v_y[0+:2],_q___pip_5160_1_91___stage___block_26_v_x[0+:2]};

_t___stage___block_1805_vnum1 = {_q___pip_5160_1_91___stage___block_26_v_z[2+:2],_q___pip_5160_1_91___stage___block_26_v_y[2+:2],_q___pip_5160_1_91___stage___block_26_v_x[2+:2]};

_t___stage___block_1805_vnum2 = {_q___pip_5160_1_91___stage___block_26_v_z[4+:2],_q___pip_5160_1_91___stage___block_26_v_y[4+:2],_q___pip_5160_1_91___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_91___stage___block_6_inside&_w_tile[_t___stage___block_1805_vnum0+:1]&_w_tile[_t___stage___block_1805_vnum1+:1]&_w_tile[_t___stage___block_1805_vnum2+:1]) begin
// __block_1806
// __block_1808
_d___pip_5160_1_91___stage___block_6_clr = _t___stage___block_1805_tex;

_d___pip_5160_1_91___stage___block_6_dist = 156;

_d___pip_5160_1_91___stage___block_6_inside = 1;

// __block_1809
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1807
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1810
_t___block_1810_cmp_yx = _q___pip_5160_1_91___block_34_tm_y-_q___pip_5160_1_91___block_34_tm_x;

_t___block_1810_cmp_zx = _q___pip_5160_1_91___block_34_tm_z-_q___pip_5160_1_91___block_34_tm_x;

_t___block_1810_cmp_zy = _q___pip_5160_1_91___block_34_tm_z-_q___pip_5160_1_91___block_34_tm_y;

_t___block_1810_x_sel = ~_t___block_1810_cmp_yx[20+:1]&&~_t___block_1810_cmp_zx[20+:1];

_t___block_1810_y_sel = _t___block_1810_cmp_yx[20+:1]&&~_t___block_1810_cmp_zy[20+:1];

_t___block_1810_z_sel = _t___block_1810_cmp_zx[20+:1]&&_t___block_1810_cmp_zy[20+:1];

if (_t___block_1810_x_sel) begin
// __block_1811
// __block_1813
_d___pip_5160_1_91___stage___block_26_v_x = _q___pip_5160_1_91___stage___block_26_v_x+_q___pip_5160_1_91___stage___block_26_s_x;

_d___pip_5160_1_91___block_34_tm_x = _q___pip_5160_1_91___block_34_tm_x+_q___pip_5160_1_91___block_40_dt_x;

// __block_1814
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1812
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1815
if (_t___block_1810_y_sel) begin
// __block_1816
// __block_1818
_d___pip_5160_1_91___stage___block_26_v_y = _q___pip_5160_1_91___stage___block_26_v_y+_q___pip_5160_1_91___stage___block_26_s_y;

_d___pip_5160_1_91___block_34_tm_y = _q___pip_5160_1_91___block_34_tm_y+_q___pip_5160_1_91___block_40_dt_y;

// __block_1819
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1817
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1820
if (_t___block_1810_z_sel) begin
// __block_1821
// __block_1823
_d___pip_5160_1_91___stage___block_26_v_z = _q___pip_5160_1_91___stage___block_26_v_z+_q___pip_5160_1_91___stage___block_26_s_z;

_d___pip_5160_1_91___block_34_tm_z = _q___pip_5160_1_91___block_34_tm_z+_q___pip_5160_1_91___block_40_dt_z;

// __block_1824
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1822
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1825
// end of pipeline stage
_d__full_fsm___pip_5160_1_91 = 1;
_d__idx_fsm___pip_5160_1_91 = _t__stall_fsm___pip_5160_1_91 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_91 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 92
(* full_case *)
case (_q__idx_fsm___pip_5160_1_92)
1: begin
// __stage___block_1826
_t___stage___block_1826_tex = (_q___pip_5160_1_92___stage___block_26_v_x)^(_q___pip_5160_1_92___stage___block_26_v_y)^(_q___pip_5160_1_92___stage___block_26_v_z);

_t___stage___block_1826_vnum0 = {_q___pip_5160_1_92___stage___block_26_v_z[0+:2],_q___pip_5160_1_92___stage___block_26_v_y[0+:2],_q___pip_5160_1_92___stage___block_26_v_x[0+:2]};

_t___stage___block_1826_vnum1 = {_q___pip_5160_1_92___stage___block_26_v_z[2+:2],_q___pip_5160_1_92___stage___block_26_v_y[2+:2],_q___pip_5160_1_92___stage___block_26_v_x[2+:2]};

_t___stage___block_1826_vnum2 = {_q___pip_5160_1_92___stage___block_26_v_z[4+:2],_q___pip_5160_1_92___stage___block_26_v_y[4+:2],_q___pip_5160_1_92___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_92___stage___block_6_inside&_w_tile[_t___stage___block_1826_vnum0+:1]&_w_tile[_t___stage___block_1826_vnum1+:1]&_w_tile[_t___stage___block_1826_vnum2+:1]) begin
// __block_1827
// __block_1829
_d___pip_5160_1_92___stage___block_6_clr = _t___stage___block_1826_tex;

_d___pip_5160_1_92___stage___block_6_dist = 158;

_d___pip_5160_1_92___stage___block_6_inside = 1;

// __block_1830
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1828
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1831
_t___block_1831_cmp_yx = _q___pip_5160_1_92___block_34_tm_y-_q___pip_5160_1_92___block_34_tm_x;

_t___block_1831_cmp_zx = _q___pip_5160_1_92___block_34_tm_z-_q___pip_5160_1_92___block_34_tm_x;

_t___block_1831_cmp_zy = _q___pip_5160_1_92___block_34_tm_z-_q___pip_5160_1_92___block_34_tm_y;

_t___block_1831_x_sel = ~_t___block_1831_cmp_yx[20+:1]&&~_t___block_1831_cmp_zx[20+:1];

_t___block_1831_y_sel = _t___block_1831_cmp_yx[20+:1]&&~_t___block_1831_cmp_zy[20+:1];

_t___block_1831_z_sel = _t___block_1831_cmp_zx[20+:1]&&_t___block_1831_cmp_zy[20+:1];

if (_t___block_1831_x_sel) begin
// __block_1832
// __block_1834
_d___pip_5160_1_92___stage___block_26_v_x = _q___pip_5160_1_92___stage___block_26_v_x+_q___pip_5160_1_92___stage___block_26_s_x;

_d___pip_5160_1_92___block_34_tm_x = _q___pip_5160_1_92___block_34_tm_x+_q___pip_5160_1_92___block_40_dt_x;

// __block_1835
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1833
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1836
if (_t___block_1831_y_sel) begin
// __block_1837
// __block_1839
_d___pip_5160_1_92___stage___block_26_v_y = _q___pip_5160_1_92___stage___block_26_v_y+_q___pip_5160_1_92___stage___block_26_s_y;

_d___pip_5160_1_92___block_34_tm_y = _q___pip_5160_1_92___block_34_tm_y+_q___pip_5160_1_92___block_40_dt_y;

// __block_1840
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1838
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1841
if (_t___block_1831_z_sel) begin
// __block_1842
// __block_1844
_d___pip_5160_1_92___stage___block_26_v_z = _q___pip_5160_1_92___stage___block_26_v_z+_q___pip_5160_1_92___stage___block_26_s_z;

_d___pip_5160_1_92___block_34_tm_z = _q___pip_5160_1_92___block_34_tm_z+_q___pip_5160_1_92___block_40_dt_z;

// __block_1845
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1843
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1846
// end of pipeline stage
_d__full_fsm___pip_5160_1_92 = 1;
_d__idx_fsm___pip_5160_1_92 = _t__stall_fsm___pip_5160_1_92 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_92 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 93
(* full_case *)
case (_q__idx_fsm___pip_5160_1_93)
1: begin
// __stage___block_1847
_t___stage___block_1847_tex = (_q___pip_5160_1_93___stage___block_26_v_x)^(_q___pip_5160_1_93___stage___block_26_v_y)^(_q___pip_5160_1_93___stage___block_26_v_z);

_t___stage___block_1847_vnum0 = {_q___pip_5160_1_93___stage___block_26_v_z[0+:2],_q___pip_5160_1_93___stage___block_26_v_y[0+:2],_q___pip_5160_1_93___stage___block_26_v_x[0+:2]};

_t___stage___block_1847_vnum1 = {_q___pip_5160_1_93___stage___block_26_v_z[2+:2],_q___pip_5160_1_93___stage___block_26_v_y[2+:2],_q___pip_5160_1_93___stage___block_26_v_x[2+:2]};

_t___stage___block_1847_vnum2 = {_q___pip_5160_1_93___stage___block_26_v_z[4+:2],_q___pip_5160_1_93___stage___block_26_v_y[4+:2],_q___pip_5160_1_93___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_93___stage___block_6_inside&_w_tile[_t___stage___block_1847_vnum0+:1]&_w_tile[_t___stage___block_1847_vnum1+:1]&_w_tile[_t___stage___block_1847_vnum2+:1]) begin
// __block_1848
// __block_1850
_d___pip_5160_1_93___stage___block_6_clr = _t___stage___block_1847_tex;

_d___pip_5160_1_93___stage___block_6_dist = 160;

_d___pip_5160_1_93___stage___block_6_inside = 1;

// __block_1851
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1849
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1852
_t___block_1852_cmp_yx = _q___pip_5160_1_93___block_34_tm_y-_q___pip_5160_1_93___block_34_tm_x;

_t___block_1852_cmp_zx = _q___pip_5160_1_93___block_34_tm_z-_q___pip_5160_1_93___block_34_tm_x;

_t___block_1852_cmp_zy = _q___pip_5160_1_93___block_34_tm_z-_q___pip_5160_1_93___block_34_tm_y;

_t___block_1852_x_sel = ~_t___block_1852_cmp_yx[20+:1]&&~_t___block_1852_cmp_zx[20+:1];

_t___block_1852_y_sel = _t___block_1852_cmp_yx[20+:1]&&~_t___block_1852_cmp_zy[20+:1];

_t___block_1852_z_sel = _t___block_1852_cmp_zx[20+:1]&&_t___block_1852_cmp_zy[20+:1];

if (_t___block_1852_x_sel) begin
// __block_1853
// __block_1855
_d___pip_5160_1_93___stage___block_26_v_x = _q___pip_5160_1_93___stage___block_26_v_x+_q___pip_5160_1_93___stage___block_26_s_x;

_d___pip_5160_1_93___block_34_tm_x = _q___pip_5160_1_93___block_34_tm_x+_q___pip_5160_1_93___block_40_dt_x;

// __block_1856
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1854
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1857
if (_t___block_1852_y_sel) begin
// __block_1858
// __block_1860
_d___pip_5160_1_93___stage___block_26_v_y = _q___pip_5160_1_93___stage___block_26_v_y+_q___pip_5160_1_93___stage___block_26_s_y;

_d___pip_5160_1_93___block_34_tm_y = _q___pip_5160_1_93___block_34_tm_y+_q___pip_5160_1_93___block_40_dt_y;

// __block_1861
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1859
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1862
if (_t___block_1852_z_sel) begin
// __block_1863
// __block_1865
_d___pip_5160_1_93___stage___block_26_v_z = _q___pip_5160_1_93___stage___block_26_v_z+_q___pip_5160_1_93___stage___block_26_s_z;

_d___pip_5160_1_93___block_34_tm_z = _q___pip_5160_1_93___block_34_tm_z+_q___pip_5160_1_93___block_40_dt_z;

// __block_1866
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1864
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1867
// end of pipeline stage
_d__full_fsm___pip_5160_1_93 = 1;
_d__idx_fsm___pip_5160_1_93 = _t__stall_fsm___pip_5160_1_93 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_93 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 94
(* full_case *)
case (_q__idx_fsm___pip_5160_1_94)
1: begin
// __stage___block_1868
_t___stage___block_1868_tex = (_q___pip_5160_1_94___stage___block_26_v_x)^(_q___pip_5160_1_94___stage___block_26_v_y)^(_q___pip_5160_1_94___stage___block_26_v_z);

_t___stage___block_1868_vnum0 = {_q___pip_5160_1_94___stage___block_26_v_z[0+:2],_q___pip_5160_1_94___stage___block_26_v_y[0+:2],_q___pip_5160_1_94___stage___block_26_v_x[0+:2]};

_t___stage___block_1868_vnum1 = {_q___pip_5160_1_94___stage___block_26_v_z[2+:2],_q___pip_5160_1_94___stage___block_26_v_y[2+:2],_q___pip_5160_1_94___stage___block_26_v_x[2+:2]};

_t___stage___block_1868_vnum2 = {_q___pip_5160_1_94___stage___block_26_v_z[4+:2],_q___pip_5160_1_94___stage___block_26_v_y[4+:2],_q___pip_5160_1_94___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_94___stage___block_6_inside&_w_tile[_t___stage___block_1868_vnum0+:1]&_w_tile[_t___stage___block_1868_vnum1+:1]&_w_tile[_t___stage___block_1868_vnum2+:1]) begin
// __block_1869
// __block_1871
_d___pip_5160_1_94___stage___block_6_clr = _t___stage___block_1868_tex;

_d___pip_5160_1_94___stage___block_6_dist = 162;

_d___pip_5160_1_94___stage___block_6_inside = 1;

// __block_1872
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1870
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1873
_t___block_1873_cmp_yx = _q___pip_5160_1_94___block_34_tm_y-_q___pip_5160_1_94___block_34_tm_x;

_t___block_1873_cmp_zx = _q___pip_5160_1_94___block_34_tm_z-_q___pip_5160_1_94___block_34_tm_x;

_t___block_1873_cmp_zy = _q___pip_5160_1_94___block_34_tm_z-_q___pip_5160_1_94___block_34_tm_y;

_t___block_1873_x_sel = ~_t___block_1873_cmp_yx[20+:1]&&~_t___block_1873_cmp_zx[20+:1];

_t___block_1873_y_sel = _t___block_1873_cmp_yx[20+:1]&&~_t___block_1873_cmp_zy[20+:1];

_t___block_1873_z_sel = _t___block_1873_cmp_zx[20+:1]&&_t___block_1873_cmp_zy[20+:1];

if (_t___block_1873_x_sel) begin
// __block_1874
// __block_1876
_d___pip_5160_1_94___stage___block_26_v_x = _q___pip_5160_1_94___stage___block_26_v_x+_q___pip_5160_1_94___stage___block_26_s_x;

_d___pip_5160_1_94___block_34_tm_x = _q___pip_5160_1_94___block_34_tm_x+_q___pip_5160_1_94___block_40_dt_x;

// __block_1877
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1875
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1878
if (_t___block_1873_y_sel) begin
// __block_1879
// __block_1881
_d___pip_5160_1_94___stage___block_26_v_y = _q___pip_5160_1_94___stage___block_26_v_y+_q___pip_5160_1_94___stage___block_26_s_y;

_d___pip_5160_1_94___block_34_tm_y = _q___pip_5160_1_94___block_34_tm_y+_q___pip_5160_1_94___block_40_dt_y;

// __block_1882
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1880
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1883
if (_t___block_1873_z_sel) begin
// __block_1884
// __block_1886
_d___pip_5160_1_94___stage___block_26_v_z = _q___pip_5160_1_94___stage___block_26_v_z+_q___pip_5160_1_94___stage___block_26_s_z;

_d___pip_5160_1_94___block_34_tm_z = _q___pip_5160_1_94___block_34_tm_z+_q___pip_5160_1_94___block_40_dt_z;

// __block_1887
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1885
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1888
// end of pipeline stage
_d__full_fsm___pip_5160_1_94 = 1;
_d__idx_fsm___pip_5160_1_94 = _t__stall_fsm___pip_5160_1_94 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_94 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 95
(* full_case *)
case (_q__idx_fsm___pip_5160_1_95)
1: begin
// __stage___block_1889
_t___stage___block_1889_tex = (_q___pip_5160_1_95___stage___block_26_v_x)^(_q___pip_5160_1_95___stage___block_26_v_y)^(_q___pip_5160_1_95___stage___block_26_v_z);

_t___stage___block_1889_vnum0 = {_q___pip_5160_1_95___stage___block_26_v_z[0+:2],_q___pip_5160_1_95___stage___block_26_v_y[0+:2],_q___pip_5160_1_95___stage___block_26_v_x[0+:2]};

_t___stage___block_1889_vnum1 = {_q___pip_5160_1_95___stage___block_26_v_z[2+:2],_q___pip_5160_1_95___stage___block_26_v_y[2+:2],_q___pip_5160_1_95___stage___block_26_v_x[2+:2]};

_t___stage___block_1889_vnum2 = {_q___pip_5160_1_95___stage___block_26_v_z[4+:2],_q___pip_5160_1_95___stage___block_26_v_y[4+:2],_q___pip_5160_1_95___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_95___stage___block_6_inside&_w_tile[_t___stage___block_1889_vnum0+:1]&_w_tile[_t___stage___block_1889_vnum1+:1]&_w_tile[_t___stage___block_1889_vnum2+:1]) begin
// __block_1890
// __block_1892
_d___pip_5160_1_95___stage___block_6_clr = _t___stage___block_1889_tex;

_d___pip_5160_1_95___stage___block_6_dist = 164;

_d___pip_5160_1_95___stage___block_6_inside = 1;

// __block_1893
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1891
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1894
_t___block_1894_cmp_yx = _q___pip_5160_1_95___block_34_tm_y-_q___pip_5160_1_95___block_34_tm_x;

_t___block_1894_cmp_zx = _q___pip_5160_1_95___block_34_tm_z-_q___pip_5160_1_95___block_34_tm_x;

_t___block_1894_cmp_zy = _q___pip_5160_1_95___block_34_tm_z-_q___pip_5160_1_95___block_34_tm_y;

_t___block_1894_x_sel = ~_t___block_1894_cmp_yx[20+:1]&&~_t___block_1894_cmp_zx[20+:1];

_t___block_1894_y_sel = _t___block_1894_cmp_yx[20+:1]&&~_t___block_1894_cmp_zy[20+:1];

_t___block_1894_z_sel = _t___block_1894_cmp_zx[20+:1]&&_t___block_1894_cmp_zy[20+:1];

if (_t___block_1894_x_sel) begin
// __block_1895
// __block_1897
_d___pip_5160_1_95___stage___block_26_v_x = _q___pip_5160_1_95___stage___block_26_v_x+_q___pip_5160_1_95___stage___block_26_s_x;

_d___pip_5160_1_95___block_34_tm_x = _q___pip_5160_1_95___block_34_tm_x+_q___pip_5160_1_95___block_40_dt_x;

// __block_1898
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1896
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1899
if (_t___block_1894_y_sel) begin
// __block_1900
// __block_1902
_d___pip_5160_1_95___stage___block_26_v_y = _q___pip_5160_1_95___stage___block_26_v_y+_q___pip_5160_1_95___stage___block_26_s_y;

_d___pip_5160_1_95___block_34_tm_y = _q___pip_5160_1_95___block_34_tm_y+_q___pip_5160_1_95___block_40_dt_y;

// __block_1903
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1901
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1904
if (_t___block_1894_z_sel) begin
// __block_1905
// __block_1907
_d___pip_5160_1_95___stage___block_26_v_z = _q___pip_5160_1_95___stage___block_26_v_z+_q___pip_5160_1_95___stage___block_26_s_z;

_d___pip_5160_1_95___block_34_tm_z = _q___pip_5160_1_95___block_34_tm_z+_q___pip_5160_1_95___block_40_dt_z;

// __block_1908
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1906
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1909
// end of pipeline stage
_d__full_fsm___pip_5160_1_95 = 1;
_d__idx_fsm___pip_5160_1_95 = _t__stall_fsm___pip_5160_1_95 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_95 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 96
(* full_case *)
case (_q__idx_fsm___pip_5160_1_96)
1: begin
// __stage___block_1910
_t___stage___block_1910_tex = (_q___pip_5160_1_96___stage___block_26_v_x)^(_q___pip_5160_1_96___stage___block_26_v_y)^(_q___pip_5160_1_96___stage___block_26_v_z);

_t___stage___block_1910_vnum0 = {_q___pip_5160_1_96___stage___block_26_v_z[0+:2],_q___pip_5160_1_96___stage___block_26_v_y[0+:2],_q___pip_5160_1_96___stage___block_26_v_x[0+:2]};

_t___stage___block_1910_vnum1 = {_q___pip_5160_1_96___stage___block_26_v_z[2+:2],_q___pip_5160_1_96___stage___block_26_v_y[2+:2],_q___pip_5160_1_96___stage___block_26_v_x[2+:2]};

_t___stage___block_1910_vnum2 = {_q___pip_5160_1_96___stage___block_26_v_z[4+:2],_q___pip_5160_1_96___stage___block_26_v_y[4+:2],_q___pip_5160_1_96___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_96___stage___block_6_inside&_w_tile[_t___stage___block_1910_vnum0+:1]&_w_tile[_t___stage___block_1910_vnum1+:1]&_w_tile[_t___stage___block_1910_vnum2+:1]) begin
// __block_1911
// __block_1913
_d___pip_5160_1_96___stage___block_6_clr = _t___stage___block_1910_tex;

_d___pip_5160_1_96___stage___block_6_dist = 166;

_d___pip_5160_1_96___stage___block_6_inside = 1;

// __block_1914
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1912
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1915
_t___block_1915_cmp_yx = _q___pip_5160_1_96___block_34_tm_y-_q___pip_5160_1_96___block_34_tm_x;

_t___block_1915_cmp_zx = _q___pip_5160_1_96___block_34_tm_z-_q___pip_5160_1_96___block_34_tm_x;

_t___block_1915_cmp_zy = _q___pip_5160_1_96___block_34_tm_z-_q___pip_5160_1_96___block_34_tm_y;

_t___block_1915_x_sel = ~_t___block_1915_cmp_yx[20+:1]&&~_t___block_1915_cmp_zx[20+:1];

_t___block_1915_y_sel = _t___block_1915_cmp_yx[20+:1]&&~_t___block_1915_cmp_zy[20+:1];

_t___block_1915_z_sel = _t___block_1915_cmp_zx[20+:1]&&_t___block_1915_cmp_zy[20+:1];

if (_t___block_1915_x_sel) begin
// __block_1916
// __block_1918
_d___pip_5160_1_96___stage___block_26_v_x = _q___pip_5160_1_96___stage___block_26_v_x+_q___pip_5160_1_96___stage___block_26_s_x;

_d___pip_5160_1_96___block_34_tm_x = _q___pip_5160_1_96___block_34_tm_x+_q___pip_5160_1_96___block_40_dt_x;

// __block_1919
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1917
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1920
if (_t___block_1915_y_sel) begin
// __block_1921
// __block_1923
_d___pip_5160_1_96___stage___block_26_v_y = _q___pip_5160_1_96___stage___block_26_v_y+_q___pip_5160_1_96___stage___block_26_s_y;

_d___pip_5160_1_96___block_34_tm_y = _q___pip_5160_1_96___block_34_tm_y+_q___pip_5160_1_96___block_40_dt_y;

// __block_1924
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1922
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1925
if (_t___block_1915_z_sel) begin
// __block_1926
// __block_1928
_d___pip_5160_1_96___stage___block_26_v_z = _q___pip_5160_1_96___stage___block_26_v_z+_q___pip_5160_1_96___stage___block_26_s_z;

_d___pip_5160_1_96___block_34_tm_z = _q___pip_5160_1_96___block_34_tm_z+_q___pip_5160_1_96___block_40_dt_z;

// __block_1929
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1927
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1930
// end of pipeline stage
_d__full_fsm___pip_5160_1_96 = 1;
_d__idx_fsm___pip_5160_1_96 = _t__stall_fsm___pip_5160_1_96 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_96 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 97
(* full_case *)
case (_q__idx_fsm___pip_5160_1_97)
1: begin
// __stage___block_1931
_t___stage___block_1931_tex = (_q___pip_5160_1_97___stage___block_26_v_x)^(_q___pip_5160_1_97___stage___block_26_v_y)^(_q___pip_5160_1_97___stage___block_26_v_z);

_t___stage___block_1931_vnum0 = {_q___pip_5160_1_97___stage___block_26_v_z[0+:2],_q___pip_5160_1_97___stage___block_26_v_y[0+:2],_q___pip_5160_1_97___stage___block_26_v_x[0+:2]};

_t___stage___block_1931_vnum1 = {_q___pip_5160_1_97___stage___block_26_v_z[2+:2],_q___pip_5160_1_97___stage___block_26_v_y[2+:2],_q___pip_5160_1_97___stage___block_26_v_x[2+:2]};

_t___stage___block_1931_vnum2 = {_q___pip_5160_1_97___stage___block_26_v_z[4+:2],_q___pip_5160_1_97___stage___block_26_v_y[4+:2],_q___pip_5160_1_97___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_97___stage___block_6_inside&_w_tile[_t___stage___block_1931_vnum0+:1]&_w_tile[_t___stage___block_1931_vnum1+:1]&_w_tile[_t___stage___block_1931_vnum2+:1]) begin
// __block_1932
// __block_1934
_d___pip_5160_1_97___stage___block_6_clr = _t___stage___block_1931_tex;

_d___pip_5160_1_97___stage___block_6_dist = 168;

_d___pip_5160_1_97___stage___block_6_inside = 1;

// __block_1935
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1933
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1936
_t___block_1936_cmp_yx = _q___pip_5160_1_97___block_34_tm_y-_q___pip_5160_1_97___block_34_tm_x;

_t___block_1936_cmp_zx = _q___pip_5160_1_97___block_34_tm_z-_q___pip_5160_1_97___block_34_tm_x;

_t___block_1936_cmp_zy = _q___pip_5160_1_97___block_34_tm_z-_q___pip_5160_1_97___block_34_tm_y;

_t___block_1936_x_sel = ~_t___block_1936_cmp_yx[20+:1]&&~_t___block_1936_cmp_zx[20+:1];

_t___block_1936_y_sel = _t___block_1936_cmp_yx[20+:1]&&~_t___block_1936_cmp_zy[20+:1];

_t___block_1936_z_sel = _t___block_1936_cmp_zx[20+:1]&&_t___block_1936_cmp_zy[20+:1];

if (_t___block_1936_x_sel) begin
// __block_1937
// __block_1939
_d___pip_5160_1_97___stage___block_26_v_x = _q___pip_5160_1_97___stage___block_26_v_x+_q___pip_5160_1_97___stage___block_26_s_x;

_d___pip_5160_1_97___block_34_tm_x = _q___pip_5160_1_97___block_34_tm_x+_q___pip_5160_1_97___block_40_dt_x;

// __block_1940
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1938
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1941
if (_t___block_1936_y_sel) begin
// __block_1942
// __block_1944
_d___pip_5160_1_97___stage___block_26_v_y = _q___pip_5160_1_97___stage___block_26_v_y+_q___pip_5160_1_97___stage___block_26_s_y;

_d___pip_5160_1_97___block_34_tm_y = _q___pip_5160_1_97___block_34_tm_y+_q___pip_5160_1_97___block_40_dt_y;

// __block_1945
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1943
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1946
if (_t___block_1936_z_sel) begin
// __block_1947
// __block_1949
_d___pip_5160_1_97___stage___block_26_v_z = _q___pip_5160_1_97___stage___block_26_v_z+_q___pip_5160_1_97___stage___block_26_s_z;

_d___pip_5160_1_97___block_34_tm_z = _q___pip_5160_1_97___block_34_tm_z+_q___pip_5160_1_97___block_40_dt_z;

// __block_1950
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1948
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1951
// end of pipeline stage
_d__full_fsm___pip_5160_1_97 = 1;
_d__idx_fsm___pip_5160_1_97 = _t__stall_fsm___pip_5160_1_97 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_97 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 98
(* full_case *)
case (_q__idx_fsm___pip_5160_1_98)
1: begin
// __stage___block_1952
_t___stage___block_1952_tex = (_q___pip_5160_1_98___stage___block_26_v_x)^(_q___pip_5160_1_98___stage___block_26_v_y)^(_q___pip_5160_1_98___stage___block_26_v_z);

_t___stage___block_1952_vnum0 = {_q___pip_5160_1_98___stage___block_26_v_z[0+:2],_q___pip_5160_1_98___stage___block_26_v_y[0+:2],_q___pip_5160_1_98___stage___block_26_v_x[0+:2]};

_t___stage___block_1952_vnum1 = {_q___pip_5160_1_98___stage___block_26_v_z[2+:2],_q___pip_5160_1_98___stage___block_26_v_y[2+:2],_q___pip_5160_1_98___stage___block_26_v_x[2+:2]};

_t___stage___block_1952_vnum2 = {_q___pip_5160_1_98___stage___block_26_v_z[4+:2],_q___pip_5160_1_98___stage___block_26_v_y[4+:2],_q___pip_5160_1_98___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_98___stage___block_6_inside&_w_tile[_t___stage___block_1952_vnum0+:1]&_w_tile[_t___stage___block_1952_vnum1+:1]&_w_tile[_t___stage___block_1952_vnum2+:1]) begin
// __block_1953
// __block_1955
_d___pip_5160_1_98___stage___block_6_clr = _t___stage___block_1952_tex;

_d___pip_5160_1_98___stage___block_6_dist = 169;

_d___pip_5160_1_98___stage___block_6_inside = 1;

// __block_1956
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1954
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1957
_t___block_1957_cmp_yx = _q___pip_5160_1_98___block_34_tm_y-_q___pip_5160_1_98___block_34_tm_x;

_t___block_1957_cmp_zx = _q___pip_5160_1_98___block_34_tm_z-_q___pip_5160_1_98___block_34_tm_x;

_t___block_1957_cmp_zy = _q___pip_5160_1_98___block_34_tm_z-_q___pip_5160_1_98___block_34_tm_y;

_t___block_1957_x_sel = ~_t___block_1957_cmp_yx[20+:1]&&~_t___block_1957_cmp_zx[20+:1];

_t___block_1957_y_sel = _t___block_1957_cmp_yx[20+:1]&&~_t___block_1957_cmp_zy[20+:1];

_t___block_1957_z_sel = _t___block_1957_cmp_zx[20+:1]&&_t___block_1957_cmp_zy[20+:1];

if (_t___block_1957_x_sel) begin
// __block_1958
// __block_1960
_d___pip_5160_1_98___stage___block_26_v_x = _q___pip_5160_1_98___stage___block_26_v_x+_q___pip_5160_1_98___stage___block_26_s_x;

_d___pip_5160_1_98___block_34_tm_x = _q___pip_5160_1_98___block_34_tm_x+_q___pip_5160_1_98___block_40_dt_x;

// __block_1961
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1959
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1962
if (_t___block_1957_y_sel) begin
// __block_1963
// __block_1965
_d___pip_5160_1_98___stage___block_26_v_y = _q___pip_5160_1_98___stage___block_26_v_y+_q___pip_5160_1_98___stage___block_26_s_y;

_d___pip_5160_1_98___block_34_tm_y = _q___pip_5160_1_98___block_34_tm_y+_q___pip_5160_1_98___block_40_dt_y;

// __block_1966
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1964
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1967
if (_t___block_1957_z_sel) begin
// __block_1968
// __block_1970
_d___pip_5160_1_98___stage___block_26_v_z = _q___pip_5160_1_98___stage___block_26_v_z+_q___pip_5160_1_98___stage___block_26_s_z;

_d___pip_5160_1_98___block_34_tm_z = _q___pip_5160_1_98___block_34_tm_z+_q___pip_5160_1_98___block_40_dt_z;

// __block_1971
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1969
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1972
// end of pipeline stage
_d__full_fsm___pip_5160_1_98 = 1;
_d__idx_fsm___pip_5160_1_98 = _t__stall_fsm___pip_5160_1_98 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_98 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 99
(* full_case *)
case (_q__idx_fsm___pip_5160_1_99)
1: begin
// __stage___block_1973
_t___stage___block_1973_tex = (_q___pip_5160_1_99___stage___block_26_v_x)^(_q___pip_5160_1_99___stage___block_26_v_y)^(_q___pip_5160_1_99___stage___block_26_v_z);

_t___stage___block_1973_vnum0 = {_q___pip_5160_1_99___stage___block_26_v_z[0+:2],_q___pip_5160_1_99___stage___block_26_v_y[0+:2],_q___pip_5160_1_99___stage___block_26_v_x[0+:2]};

_t___stage___block_1973_vnum1 = {_q___pip_5160_1_99___stage___block_26_v_z[2+:2],_q___pip_5160_1_99___stage___block_26_v_y[2+:2],_q___pip_5160_1_99___stage___block_26_v_x[2+:2]};

_t___stage___block_1973_vnum2 = {_q___pip_5160_1_99___stage___block_26_v_z[4+:2],_q___pip_5160_1_99___stage___block_26_v_y[4+:2],_q___pip_5160_1_99___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_99___stage___block_6_inside&_w_tile[_t___stage___block_1973_vnum0+:1]&_w_tile[_t___stage___block_1973_vnum1+:1]&_w_tile[_t___stage___block_1973_vnum2+:1]) begin
// __block_1974
// __block_1976
_d___pip_5160_1_99___stage___block_6_clr = _t___stage___block_1973_tex;

_d___pip_5160_1_99___stage___block_6_dist = 171;

_d___pip_5160_1_99___stage___block_6_inside = 1;

// __block_1977
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1975
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1978
_t___block_1978_cmp_yx = _q___pip_5160_1_99___block_34_tm_y-_q___pip_5160_1_99___block_34_tm_x;

_t___block_1978_cmp_zx = _q___pip_5160_1_99___block_34_tm_z-_q___pip_5160_1_99___block_34_tm_x;

_t___block_1978_cmp_zy = _q___pip_5160_1_99___block_34_tm_z-_q___pip_5160_1_99___block_34_tm_y;

_t___block_1978_x_sel = ~_t___block_1978_cmp_yx[20+:1]&&~_t___block_1978_cmp_zx[20+:1];

_t___block_1978_y_sel = _t___block_1978_cmp_yx[20+:1]&&~_t___block_1978_cmp_zy[20+:1];

_t___block_1978_z_sel = _t___block_1978_cmp_zx[20+:1]&&_t___block_1978_cmp_zy[20+:1];

if (_t___block_1978_x_sel) begin
// __block_1979
// __block_1981
_d___pip_5160_1_99___stage___block_26_v_x = _q___pip_5160_1_99___stage___block_26_v_x+_q___pip_5160_1_99___stage___block_26_s_x;

_d___pip_5160_1_99___block_34_tm_x = _q___pip_5160_1_99___block_34_tm_x+_q___pip_5160_1_99___block_40_dt_x;

// __block_1982
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1980
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1983
if (_t___block_1978_y_sel) begin
// __block_1984
// __block_1986
_d___pip_5160_1_99___stage___block_26_v_y = _q___pip_5160_1_99___stage___block_26_v_y+_q___pip_5160_1_99___stage___block_26_s_y;

_d___pip_5160_1_99___block_34_tm_y = _q___pip_5160_1_99___block_34_tm_y+_q___pip_5160_1_99___block_40_dt_y;

// __block_1987
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1985
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1988
if (_t___block_1978_z_sel) begin
// __block_1989
// __block_1991
_d___pip_5160_1_99___stage___block_26_v_z = _q___pip_5160_1_99___stage___block_26_v_z+_q___pip_5160_1_99___stage___block_26_s_z;

_d___pip_5160_1_99___block_34_tm_z = _q___pip_5160_1_99___block_34_tm_z+_q___pip_5160_1_99___block_40_dt_z;

// __block_1992
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1990
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1993
// end of pipeline stage
_d__full_fsm___pip_5160_1_99 = 1;
_d__idx_fsm___pip_5160_1_99 = _t__stall_fsm___pip_5160_1_99 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_99 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 100
(* full_case *)
case (_q__idx_fsm___pip_5160_1_100)
1: begin
// __stage___block_1994
_t___stage___block_1994_tex = (_q___pip_5160_1_100___stage___block_26_v_x)^(_q___pip_5160_1_100___stage___block_26_v_y)^(_q___pip_5160_1_100___stage___block_26_v_z);

_t___stage___block_1994_vnum0 = {_q___pip_5160_1_100___stage___block_26_v_z[0+:2],_q___pip_5160_1_100___stage___block_26_v_y[0+:2],_q___pip_5160_1_100___stage___block_26_v_x[0+:2]};

_t___stage___block_1994_vnum1 = {_q___pip_5160_1_100___stage___block_26_v_z[2+:2],_q___pip_5160_1_100___stage___block_26_v_y[2+:2],_q___pip_5160_1_100___stage___block_26_v_x[2+:2]};

_t___stage___block_1994_vnum2 = {_q___pip_5160_1_100___stage___block_26_v_z[4+:2],_q___pip_5160_1_100___stage___block_26_v_y[4+:2],_q___pip_5160_1_100___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_100___stage___block_6_inside&_w_tile[_t___stage___block_1994_vnum0+:1]&_w_tile[_t___stage___block_1994_vnum1+:1]&_w_tile[_t___stage___block_1994_vnum2+:1]) begin
// __block_1995
// __block_1997
_d___pip_5160_1_100___stage___block_6_clr = _t___stage___block_1994_tex;

_d___pip_5160_1_100___stage___block_6_dist = 173;

_d___pip_5160_1_100___stage___block_6_inside = 1;

// __block_1998
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_1996
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_1999
_t___block_1999_cmp_yx = _q___pip_5160_1_100___block_34_tm_y-_q___pip_5160_1_100___block_34_tm_x;

_t___block_1999_cmp_zx = _q___pip_5160_1_100___block_34_tm_z-_q___pip_5160_1_100___block_34_tm_x;

_t___block_1999_cmp_zy = _q___pip_5160_1_100___block_34_tm_z-_q___pip_5160_1_100___block_34_tm_y;

_t___block_1999_x_sel = ~_t___block_1999_cmp_yx[20+:1]&&~_t___block_1999_cmp_zx[20+:1];

_t___block_1999_y_sel = _t___block_1999_cmp_yx[20+:1]&&~_t___block_1999_cmp_zy[20+:1];

_t___block_1999_z_sel = _t___block_1999_cmp_zx[20+:1]&&_t___block_1999_cmp_zy[20+:1];

if (_t___block_1999_x_sel) begin
// __block_2000
// __block_2002
_d___pip_5160_1_100___stage___block_26_v_x = _q___pip_5160_1_100___stage___block_26_v_x+_q___pip_5160_1_100___stage___block_26_s_x;

_d___pip_5160_1_100___block_34_tm_x = _q___pip_5160_1_100___block_34_tm_x+_q___pip_5160_1_100___block_40_dt_x;

// __block_2003
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2001
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2004
if (_t___block_1999_y_sel) begin
// __block_2005
// __block_2007
_d___pip_5160_1_100___stage___block_26_v_y = _q___pip_5160_1_100___stage___block_26_v_y+_q___pip_5160_1_100___stage___block_26_s_y;

_d___pip_5160_1_100___block_34_tm_y = _q___pip_5160_1_100___block_34_tm_y+_q___pip_5160_1_100___block_40_dt_y;

// __block_2008
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2006
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2009
if (_t___block_1999_z_sel) begin
// __block_2010
// __block_2012
_d___pip_5160_1_100___stage___block_26_v_z = _q___pip_5160_1_100___stage___block_26_v_z+_q___pip_5160_1_100___stage___block_26_s_z;

_d___pip_5160_1_100___block_34_tm_z = _q___pip_5160_1_100___block_34_tm_z+_q___pip_5160_1_100___block_40_dt_z;

// __block_2013
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2011
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2014
// end of pipeline stage
_d__full_fsm___pip_5160_1_100 = 1;
_d__idx_fsm___pip_5160_1_100 = _t__stall_fsm___pip_5160_1_100 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_100 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 101
(* full_case *)
case (_q__idx_fsm___pip_5160_1_101)
1: begin
// __stage___block_2015
_t___stage___block_2015_tex = (_q___pip_5160_1_101___stage___block_26_v_x)^(_q___pip_5160_1_101___stage___block_26_v_y)^(_q___pip_5160_1_101___stage___block_26_v_z);

_t___stage___block_2015_vnum0 = {_q___pip_5160_1_101___stage___block_26_v_z[0+:2],_q___pip_5160_1_101___stage___block_26_v_y[0+:2],_q___pip_5160_1_101___stage___block_26_v_x[0+:2]};

_t___stage___block_2015_vnum1 = {_q___pip_5160_1_101___stage___block_26_v_z[2+:2],_q___pip_5160_1_101___stage___block_26_v_y[2+:2],_q___pip_5160_1_101___stage___block_26_v_x[2+:2]};

_t___stage___block_2015_vnum2 = {_q___pip_5160_1_101___stage___block_26_v_z[4+:2],_q___pip_5160_1_101___stage___block_26_v_y[4+:2],_q___pip_5160_1_101___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_101___stage___block_6_inside&_w_tile[_t___stage___block_2015_vnum0+:1]&_w_tile[_t___stage___block_2015_vnum1+:1]&_w_tile[_t___stage___block_2015_vnum2+:1]) begin
// __block_2016
// __block_2018
_d___pip_5160_1_101___stage___block_6_clr = _t___stage___block_2015_tex;

_d___pip_5160_1_101___stage___block_6_dist = 175;

_d___pip_5160_1_101___stage___block_6_inside = 1;

// __block_2019
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2017
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2020
_t___block_2020_cmp_yx = _q___pip_5160_1_101___block_34_tm_y-_q___pip_5160_1_101___block_34_tm_x;

_t___block_2020_cmp_zx = _q___pip_5160_1_101___block_34_tm_z-_q___pip_5160_1_101___block_34_tm_x;

_t___block_2020_cmp_zy = _q___pip_5160_1_101___block_34_tm_z-_q___pip_5160_1_101___block_34_tm_y;

_t___block_2020_x_sel = ~_t___block_2020_cmp_yx[20+:1]&&~_t___block_2020_cmp_zx[20+:1];

_t___block_2020_y_sel = _t___block_2020_cmp_yx[20+:1]&&~_t___block_2020_cmp_zy[20+:1];

_t___block_2020_z_sel = _t___block_2020_cmp_zx[20+:1]&&_t___block_2020_cmp_zy[20+:1];

if (_t___block_2020_x_sel) begin
// __block_2021
// __block_2023
_d___pip_5160_1_101___stage___block_26_v_x = _q___pip_5160_1_101___stage___block_26_v_x+_q___pip_5160_1_101___stage___block_26_s_x;

_d___pip_5160_1_101___block_34_tm_x = _q___pip_5160_1_101___block_34_tm_x+_q___pip_5160_1_101___block_40_dt_x;

// __block_2024
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2022
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2025
if (_t___block_2020_y_sel) begin
// __block_2026
// __block_2028
_d___pip_5160_1_101___stage___block_26_v_y = _q___pip_5160_1_101___stage___block_26_v_y+_q___pip_5160_1_101___stage___block_26_s_y;

_d___pip_5160_1_101___block_34_tm_y = _q___pip_5160_1_101___block_34_tm_y+_q___pip_5160_1_101___block_40_dt_y;

// __block_2029
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2027
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2030
if (_t___block_2020_z_sel) begin
// __block_2031
// __block_2033
_d___pip_5160_1_101___stage___block_26_v_z = _q___pip_5160_1_101___stage___block_26_v_z+_q___pip_5160_1_101___stage___block_26_s_z;

_d___pip_5160_1_101___block_34_tm_z = _q___pip_5160_1_101___block_34_tm_z+_q___pip_5160_1_101___block_40_dt_z;

// __block_2034
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2032
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2035
// end of pipeline stage
_d__full_fsm___pip_5160_1_101 = 1;
_d__idx_fsm___pip_5160_1_101 = _t__stall_fsm___pip_5160_1_101 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_101 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 102
(* full_case *)
case (_q__idx_fsm___pip_5160_1_102)
1: begin
// __stage___block_2036
_t___stage___block_2036_tex = (_q___pip_5160_1_102___stage___block_26_v_x)^(_q___pip_5160_1_102___stage___block_26_v_y)^(_q___pip_5160_1_102___stage___block_26_v_z);

_t___stage___block_2036_vnum0 = {_q___pip_5160_1_102___stage___block_26_v_z[0+:2],_q___pip_5160_1_102___stage___block_26_v_y[0+:2],_q___pip_5160_1_102___stage___block_26_v_x[0+:2]};

_t___stage___block_2036_vnum1 = {_q___pip_5160_1_102___stage___block_26_v_z[2+:2],_q___pip_5160_1_102___stage___block_26_v_y[2+:2],_q___pip_5160_1_102___stage___block_26_v_x[2+:2]};

_t___stage___block_2036_vnum2 = {_q___pip_5160_1_102___stage___block_26_v_z[4+:2],_q___pip_5160_1_102___stage___block_26_v_y[4+:2],_q___pip_5160_1_102___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_102___stage___block_6_inside&_w_tile[_t___stage___block_2036_vnum0+:1]&_w_tile[_t___stage___block_2036_vnum1+:1]&_w_tile[_t___stage___block_2036_vnum2+:1]) begin
// __block_2037
// __block_2039
_d___pip_5160_1_102___stage___block_6_clr = _t___stage___block_2036_tex;

_d___pip_5160_1_102___stage___block_6_dist = 177;

_d___pip_5160_1_102___stage___block_6_inside = 1;

// __block_2040
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2038
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2041
_t___block_2041_cmp_yx = _q___pip_5160_1_102___block_34_tm_y-_q___pip_5160_1_102___block_34_tm_x;

_t___block_2041_cmp_zx = _q___pip_5160_1_102___block_34_tm_z-_q___pip_5160_1_102___block_34_tm_x;

_t___block_2041_cmp_zy = _q___pip_5160_1_102___block_34_tm_z-_q___pip_5160_1_102___block_34_tm_y;

_t___block_2041_x_sel = ~_t___block_2041_cmp_yx[20+:1]&&~_t___block_2041_cmp_zx[20+:1];

_t___block_2041_y_sel = _t___block_2041_cmp_yx[20+:1]&&~_t___block_2041_cmp_zy[20+:1];

_t___block_2041_z_sel = _t___block_2041_cmp_zx[20+:1]&&_t___block_2041_cmp_zy[20+:1];

if (_t___block_2041_x_sel) begin
// __block_2042
// __block_2044
_d___pip_5160_1_102___stage___block_26_v_x = _q___pip_5160_1_102___stage___block_26_v_x+_q___pip_5160_1_102___stage___block_26_s_x;

_d___pip_5160_1_102___block_34_tm_x = _q___pip_5160_1_102___block_34_tm_x+_q___pip_5160_1_102___block_40_dt_x;

// __block_2045
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2043
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2046
if (_t___block_2041_y_sel) begin
// __block_2047
// __block_2049
_d___pip_5160_1_102___stage___block_26_v_y = _q___pip_5160_1_102___stage___block_26_v_y+_q___pip_5160_1_102___stage___block_26_s_y;

_d___pip_5160_1_102___block_34_tm_y = _q___pip_5160_1_102___block_34_tm_y+_q___pip_5160_1_102___block_40_dt_y;

// __block_2050
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2048
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2051
if (_t___block_2041_z_sel) begin
// __block_2052
// __block_2054
_d___pip_5160_1_102___stage___block_26_v_z = _q___pip_5160_1_102___stage___block_26_v_z+_q___pip_5160_1_102___stage___block_26_s_z;

_d___pip_5160_1_102___block_34_tm_z = _q___pip_5160_1_102___block_34_tm_z+_q___pip_5160_1_102___block_40_dt_z;

// __block_2055
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2053
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2056
// end of pipeline stage
_d__full_fsm___pip_5160_1_102 = 1;
_d__idx_fsm___pip_5160_1_102 = _t__stall_fsm___pip_5160_1_102 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_102 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 103
(* full_case *)
case (_q__idx_fsm___pip_5160_1_103)
1: begin
// __stage___block_2057
_t___stage___block_2057_tex = (_q___pip_5160_1_103___stage___block_26_v_x)^(_q___pip_5160_1_103___stage___block_26_v_y)^(_q___pip_5160_1_103___stage___block_26_v_z);

_t___stage___block_2057_vnum0 = {_q___pip_5160_1_103___stage___block_26_v_z[0+:2],_q___pip_5160_1_103___stage___block_26_v_y[0+:2],_q___pip_5160_1_103___stage___block_26_v_x[0+:2]};

_t___stage___block_2057_vnum1 = {_q___pip_5160_1_103___stage___block_26_v_z[2+:2],_q___pip_5160_1_103___stage___block_26_v_y[2+:2],_q___pip_5160_1_103___stage___block_26_v_x[2+:2]};

_t___stage___block_2057_vnum2 = {_q___pip_5160_1_103___stage___block_26_v_z[4+:2],_q___pip_5160_1_103___stage___block_26_v_y[4+:2],_q___pip_5160_1_103___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_103___stage___block_6_inside&_w_tile[_t___stage___block_2057_vnum0+:1]&_w_tile[_t___stage___block_2057_vnum1+:1]&_w_tile[_t___stage___block_2057_vnum2+:1]) begin
// __block_2058
// __block_2060
_d___pip_5160_1_103___stage___block_6_clr = _t___stage___block_2057_tex;

_d___pip_5160_1_103___stage___block_6_dist = 179;

_d___pip_5160_1_103___stage___block_6_inside = 1;

// __block_2061
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2059
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2062
_t___block_2062_cmp_yx = _q___pip_5160_1_103___block_34_tm_y-_q___pip_5160_1_103___block_34_tm_x;

_t___block_2062_cmp_zx = _q___pip_5160_1_103___block_34_tm_z-_q___pip_5160_1_103___block_34_tm_x;

_t___block_2062_cmp_zy = _q___pip_5160_1_103___block_34_tm_z-_q___pip_5160_1_103___block_34_tm_y;

_t___block_2062_x_sel = ~_t___block_2062_cmp_yx[20+:1]&&~_t___block_2062_cmp_zx[20+:1];

_t___block_2062_y_sel = _t___block_2062_cmp_yx[20+:1]&&~_t___block_2062_cmp_zy[20+:1];

_t___block_2062_z_sel = _t___block_2062_cmp_zx[20+:1]&&_t___block_2062_cmp_zy[20+:1];

if (_t___block_2062_x_sel) begin
// __block_2063
// __block_2065
_d___pip_5160_1_103___stage___block_26_v_x = _q___pip_5160_1_103___stage___block_26_v_x+_q___pip_5160_1_103___stage___block_26_s_x;

_d___pip_5160_1_103___block_34_tm_x = _q___pip_5160_1_103___block_34_tm_x+_q___pip_5160_1_103___block_40_dt_x;

// __block_2066
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2064
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2067
if (_t___block_2062_y_sel) begin
// __block_2068
// __block_2070
_d___pip_5160_1_103___stage___block_26_v_y = _q___pip_5160_1_103___stage___block_26_v_y+_q___pip_5160_1_103___stage___block_26_s_y;

_d___pip_5160_1_103___block_34_tm_y = _q___pip_5160_1_103___block_34_tm_y+_q___pip_5160_1_103___block_40_dt_y;

// __block_2071
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2069
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2072
if (_t___block_2062_z_sel) begin
// __block_2073
// __block_2075
_d___pip_5160_1_103___stage___block_26_v_z = _q___pip_5160_1_103___stage___block_26_v_z+_q___pip_5160_1_103___stage___block_26_s_z;

_d___pip_5160_1_103___block_34_tm_z = _q___pip_5160_1_103___block_34_tm_z+_q___pip_5160_1_103___block_40_dt_z;

// __block_2076
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2074
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2077
// end of pipeline stage
_d__full_fsm___pip_5160_1_103 = 1;
_d__idx_fsm___pip_5160_1_103 = _t__stall_fsm___pip_5160_1_103 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_103 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 104
(* full_case *)
case (_q__idx_fsm___pip_5160_1_104)
1: begin
// __stage___block_2078
_t___stage___block_2078_tex = (_q___pip_5160_1_104___stage___block_26_v_x)^(_q___pip_5160_1_104___stage___block_26_v_y)^(_q___pip_5160_1_104___stage___block_26_v_z);

_t___stage___block_2078_vnum0 = {_q___pip_5160_1_104___stage___block_26_v_z[0+:2],_q___pip_5160_1_104___stage___block_26_v_y[0+:2],_q___pip_5160_1_104___stage___block_26_v_x[0+:2]};

_t___stage___block_2078_vnum1 = {_q___pip_5160_1_104___stage___block_26_v_z[2+:2],_q___pip_5160_1_104___stage___block_26_v_y[2+:2],_q___pip_5160_1_104___stage___block_26_v_x[2+:2]};

_t___stage___block_2078_vnum2 = {_q___pip_5160_1_104___stage___block_26_v_z[4+:2],_q___pip_5160_1_104___stage___block_26_v_y[4+:2],_q___pip_5160_1_104___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_104___stage___block_6_inside&_w_tile[_t___stage___block_2078_vnum0+:1]&_w_tile[_t___stage___block_2078_vnum1+:1]&_w_tile[_t___stage___block_2078_vnum2+:1]) begin
// __block_2079
// __block_2081
_d___pip_5160_1_104___stage___block_6_clr = _t___stage___block_2078_tex;

_d___pip_5160_1_104___stage___block_6_dist = 181;

_d___pip_5160_1_104___stage___block_6_inside = 1;

// __block_2082
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2080
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2083
_t___block_2083_cmp_yx = _q___pip_5160_1_104___block_34_tm_y-_q___pip_5160_1_104___block_34_tm_x;

_t___block_2083_cmp_zx = _q___pip_5160_1_104___block_34_tm_z-_q___pip_5160_1_104___block_34_tm_x;

_t___block_2083_cmp_zy = _q___pip_5160_1_104___block_34_tm_z-_q___pip_5160_1_104___block_34_tm_y;

_t___block_2083_x_sel = ~_t___block_2083_cmp_yx[20+:1]&&~_t___block_2083_cmp_zx[20+:1];

_t___block_2083_y_sel = _t___block_2083_cmp_yx[20+:1]&&~_t___block_2083_cmp_zy[20+:1];

_t___block_2083_z_sel = _t___block_2083_cmp_zx[20+:1]&&_t___block_2083_cmp_zy[20+:1];

if (_t___block_2083_x_sel) begin
// __block_2084
// __block_2086
_d___pip_5160_1_104___stage___block_26_v_x = _q___pip_5160_1_104___stage___block_26_v_x+_q___pip_5160_1_104___stage___block_26_s_x;

_d___pip_5160_1_104___block_34_tm_x = _q___pip_5160_1_104___block_34_tm_x+_q___pip_5160_1_104___block_40_dt_x;

// __block_2087
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2085
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2088
if (_t___block_2083_y_sel) begin
// __block_2089
// __block_2091
_d___pip_5160_1_104___stage___block_26_v_y = _q___pip_5160_1_104___stage___block_26_v_y+_q___pip_5160_1_104___stage___block_26_s_y;

_d___pip_5160_1_104___block_34_tm_y = _q___pip_5160_1_104___block_34_tm_y+_q___pip_5160_1_104___block_40_dt_y;

// __block_2092
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2090
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2093
if (_t___block_2083_z_sel) begin
// __block_2094
// __block_2096
_d___pip_5160_1_104___stage___block_26_v_z = _q___pip_5160_1_104___stage___block_26_v_z+_q___pip_5160_1_104___stage___block_26_s_z;

_d___pip_5160_1_104___block_34_tm_z = _q___pip_5160_1_104___block_34_tm_z+_q___pip_5160_1_104___block_40_dt_z;

// __block_2097
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2095
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2098
// end of pipeline stage
_d__full_fsm___pip_5160_1_104 = 1;
_d__idx_fsm___pip_5160_1_104 = _t__stall_fsm___pip_5160_1_104 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_104 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 105
(* full_case *)
case (_q__idx_fsm___pip_5160_1_105)
1: begin
// __stage___block_2099
_t___stage___block_2099_tex = (_q___pip_5160_1_105___stage___block_26_v_x)^(_q___pip_5160_1_105___stage___block_26_v_y)^(_q___pip_5160_1_105___stage___block_26_v_z);

_t___stage___block_2099_vnum0 = {_q___pip_5160_1_105___stage___block_26_v_z[0+:2],_q___pip_5160_1_105___stage___block_26_v_y[0+:2],_q___pip_5160_1_105___stage___block_26_v_x[0+:2]};

_t___stage___block_2099_vnum1 = {_q___pip_5160_1_105___stage___block_26_v_z[2+:2],_q___pip_5160_1_105___stage___block_26_v_y[2+:2],_q___pip_5160_1_105___stage___block_26_v_x[2+:2]};

_t___stage___block_2099_vnum2 = {_q___pip_5160_1_105___stage___block_26_v_z[4+:2],_q___pip_5160_1_105___stage___block_26_v_y[4+:2],_q___pip_5160_1_105___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_105___stage___block_6_inside&_w_tile[_t___stage___block_2099_vnum0+:1]&_w_tile[_t___stage___block_2099_vnum1+:1]&_w_tile[_t___stage___block_2099_vnum2+:1]) begin
// __block_2100
// __block_2102
_d___pip_5160_1_105___stage___block_6_clr = _t___stage___block_2099_tex;

_d___pip_5160_1_105___stage___block_6_dist = 182;

_d___pip_5160_1_105___stage___block_6_inside = 1;

// __block_2103
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2101
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2104
_t___block_2104_cmp_yx = _q___pip_5160_1_105___block_34_tm_y-_q___pip_5160_1_105___block_34_tm_x;

_t___block_2104_cmp_zx = _q___pip_5160_1_105___block_34_tm_z-_q___pip_5160_1_105___block_34_tm_x;

_t___block_2104_cmp_zy = _q___pip_5160_1_105___block_34_tm_z-_q___pip_5160_1_105___block_34_tm_y;

_t___block_2104_x_sel = ~_t___block_2104_cmp_yx[20+:1]&&~_t___block_2104_cmp_zx[20+:1];

_t___block_2104_y_sel = _t___block_2104_cmp_yx[20+:1]&&~_t___block_2104_cmp_zy[20+:1];

_t___block_2104_z_sel = _t___block_2104_cmp_zx[20+:1]&&_t___block_2104_cmp_zy[20+:1];

if (_t___block_2104_x_sel) begin
// __block_2105
// __block_2107
_d___pip_5160_1_105___stage___block_26_v_x = _q___pip_5160_1_105___stage___block_26_v_x+_q___pip_5160_1_105___stage___block_26_s_x;

_d___pip_5160_1_105___block_34_tm_x = _q___pip_5160_1_105___block_34_tm_x+_q___pip_5160_1_105___block_40_dt_x;

// __block_2108
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2106
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2109
if (_t___block_2104_y_sel) begin
// __block_2110
// __block_2112
_d___pip_5160_1_105___stage___block_26_v_y = _q___pip_5160_1_105___stage___block_26_v_y+_q___pip_5160_1_105___stage___block_26_s_y;

_d___pip_5160_1_105___block_34_tm_y = _q___pip_5160_1_105___block_34_tm_y+_q___pip_5160_1_105___block_40_dt_y;

// __block_2113
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2111
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2114
if (_t___block_2104_z_sel) begin
// __block_2115
// __block_2117
_d___pip_5160_1_105___stage___block_26_v_z = _q___pip_5160_1_105___stage___block_26_v_z+_q___pip_5160_1_105___stage___block_26_s_z;

_d___pip_5160_1_105___block_34_tm_z = _q___pip_5160_1_105___block_34_tm_z+_q___pip_5160_1_105___block_40_dt_z;

// __block_2118
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2116
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2119
// end of pipeline stage
_d__full_fsm___pip_5160_1_105 = 1;
_d__idx_fsm___pip_5160_1_105 = _t__stall_fsm___pip_5160_1_105 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_105 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 106
(* full_case *)
case (_q__idx_fsm___pip_5160_1_106)
1: begin
// __stage___block_2120
_t___stage___block_2120_tex = (_q___pip_5160_1_106___stage___block_26_v_x)^(_q___pip_5160_1_106___stage___block_26_v_y)^(_q___pip_5160_1_106___stage___block_26_v_z);

_t___stage___block_2120_vnum0 = {_q___pip_5160_1_106___stage___block_26_v_z[0+:2],_q___pip_5160_1_106___stage___block_26_v_y[0+:2],_q___pip_5160_1_106___stage___block_26_v_x[0+:2]};

_t___stage___block_2120_vnum1 = {_q___pip_5160_1_106___stage___block_26_v_z[2+:2],_q___pip_5160_1_106___stage___block_26_v_y[2+:2],_q___pip_5160_1_106___stage___block_26_v_x[2+:2]};

_t___stage___block_2120_vnum2 = {_q___pip_5160_1_106___stage___block_26_v_z[4+:2],_q___pip_5160_1_106___stage___block_26_v_y[4+:2],_q___pip_5160_1_106___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_106___stage___block_6_inside&_w_tile[_t___stage___block_2120_vnum0+:1]&_w_tile[_t___stage___block_2120_vnum1+:1]&_w_tile[_t___stage___block_2120_vnum2+:1]) begin
// __block_2121
// __block_2123
_d___pip_5160_1_106___stage___block_6_clr = _t___stage___block_2120_tex;

_d___pip_5160_1_106___stage___block_6_dist = 184;

_d___pip_5160_1_106___stage___block_6_inside = 1;

// __block_2124
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2122
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2125
_t___block_2125_cmp_yx = _q___pip_5160_1_106___block_34_tm_y-_q___pip_5160_1_106___block_34_tm_x;

_t___block_2125_cmp_zx = _q___pip_5160_1_106___block_34_tm_z-_q___pip_5160_1_106___block_34_tm_x;

_t___block_2125_cmp_zy = _q___pip_5160_1_106___block_34_tm_z-_q___pip_5160_1_106___block_34_tm_y;

_t___block_2125_x_sel = ~_t___block_2125_cmp_yx[20+:1]&&~_t___block_2125_cmp_zx[20+:1];

_t___block_2125_y_sel = _t___block_2125_cmp_yx[20+:1]&&~_t___block_2125_cmp_zy[20+:1];

_t___block_2125_z_sel = _t___block_2125_cmp_zx[20+:1]&&_t___block_2125_cmp_zy[20+:1];

if (_t___block_2125_x_sel) begin
// __block_2126
// __block_2128
_d___pip_5160_1_106___stage___block_26_v_x = _q___pip_5160_1_106___stage___block_26_v_x+_q___pip_5160_1_106___stage___block_26_s_x;

_d___pip_5160_1_106___block_34_tm_x = _q___pip_5160_1_106___block_34_tm_x+_q___pip_5160_1_106___block_40_dt_x;

// __block_2129
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2127
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2130
if (_t___block_2125_y_sel) begin
// __block_2131
// __block_2133
_d___pip_5160_1_106___stage___block_26_v_y = _q___pip_5160_1_106___stage___block_26_v_y+_q___pip_5160_1_106___stage___block_26_s_y;

_d___pip_5160_1_106___block_34_tm_y = _q___pip_5160_1_106___block_34_tm_y+_q___pip_5160_1_106___block_40_dt_y;

// __block_2134
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2132
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2135
if (_t___block_2125_z_sel) begin
// __block_2136
// __block_2138
_d___pip_5160_1_106___stage___block_26_v_z = _q___pip_5160_1_106___stage___block_26_v_z+_q___pip_5160_1_106___stage___block_26_s_z;

_d___pip_5160_1_106___block_34_tm_z = _q___pip_5160_1_106___block_34_tm_z+_q___pip_5160_1_106___block_40_dt_z;

// __block_2139
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2137
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2140
// end of pipeline stage
_d__full_fsm___pip_5160_1_106 = 1;
_d__idx_fsm___pip_5160_1_106 = _t__stall_fsm___pip_5160_1_106 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_106 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 107
(* full_case *)
case (_q__idx_fsm___pip_5160_1_107)
1: begin
// __stage___block_2141
_t___stage___block_2141_tex = (_q___pip_5160_1_107___stage___block_26_v_x)^(_q___pip_5160_1_107___stage___block_26_v_y)^(_q___pip_5160_1_107___stage___block_26_v_z);

_t___stage___block_2141_vnum0 = {_q___pip_5160_1_107___stage___block_26_v_z[0+:2],_q___pip_5160_1_107___stage___block_26_v_y[0+:2],_q___pip_5160_1_107___stage___block_26_v_x[0+:2]};

_t___stage___block_2141_vnum1 = {_q___pip_5160_1_107___stage___block_26_v_z[2+:2],_q___pip_5160_1_107___stage___block_26_v_y[2+:2],_q___pip_5160_1_107___stage___block_26_v_x[2+:2]};

_t___stage___block_2141_vnum2 = {_q___pip_5160_1_107___stage___block_26_v_z[4+:2],_q___pip_5160_1_107___stage___block_26_v_y[4+:2],_q___pip_5160_1_107___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_107___stage___block_6_inside&_w_tile[_t___stage___block_2141_vnum0+:1]&_w_tile[_t___stage___block_2141_vnum1+:1]&_w_tile[_t___stage___block_2141_vnum2+:1]) begin
// __block_2142
// __block_2144
_d___pip_5160_1_107___stage___block_6_clr = _t___stage___block_2141_tex;

_d___pip_5160_1_107___stage___block_6_dist = 186;

_d___pip_5160_1_107___stage___block_6_inside = 1;

// __block_2145
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2143
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2146
_t___block_2146_cmp_yx = _q___pip_5160_1_107___block_34_tm_y-_q___pip_5160_1_107___block_34_tm_x;

_t___block_2146_cmp_zx = _q___pip_5160_1_107___block_34_tm_z-_q___pip_5160_1_107___block_34_tm_x;

_t___block_2146_cmp_zy = _q___pip_5160_1_107___block_34_tm_z-_q___pip_5160_1_107___block_34_tm_y;

_t___block_2146_x_sel = ~_t___block_2146_cmp_yx[20+:1]&&~_t___block_2146_cmp_zx[20+:1];

_t___block_2146_y_sel = _t___block_2146_cmp_yx[20+:1]&&~_t___block_2146_cmp_zy[20+:1];

_t___block_2146_z_sel = _t___block_2146_cmp_zx[20+:1]&&_t___block_2146_cmp_zy[20+:1];

if (_t___block_2146_x_sel) begin
// __block_2147
// __block_2149
_d___pip_5160_1_107___stage___block_26_v_x = _q___pip_5160_1_107___stage___block_26_v_x+_q___pip_5160_1_107___stage___block_26_s_x;

_d___pip_5160_1_107___block_34_tm_x = _q___pip_5160_1_107___block_34_tm_x+_q___pip_5160_1_107___block_40_dt_x;

// __block_2150
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2148
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2151
if (_t___block_2146_y_sel) begin
// __block_2152
// __block_2154
_d___pip_5160_1_107___stage___block_26_v_y = _q___pip_5160_1_107___stage___block_26_v_y+_q___pip_5160_1_107___stage___block_26_s_y;

_d___pip_5160_1_107___block_34_tm_y = _q___pip_5160_1_107___block_34_tm_y+_q___pip_5160_1_107___block_40_dt_y;

// __block_2155
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2153
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2156
if (_t___block_2146_z_sel) begin
// __block_2157
// __block_2159
_d___pip_5160_1_107___stage___block_26_v_z = _q___pip_5160_1_107___stage___block_26_v_z+_q___pip_5160_1_107___stage___block_26_s_z;

_d___pip_5160_1_107___block_34_tm_z = _q___pip_5160_1_107___block_34_tm_z+_q___pip_5160_1_107___block_40_dt_z;

// __block_2160
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2158
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2161
// end of pipeline stage
_d__full_fsm___pip_5160_1_107 = 1;
_d__idx_fsm___pip_5160_1_107 = _t__stall_fsm___pip_5160_1_107 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_107 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 108
(* full_case *)
case (_q__idx_fsm___pip_5160_1_108)
1: begin
// __stage___block_2162
_t___stage___block_2162_tex = (_q___pip_5160_1_108___stage___block_26_v_x)^(_q___pip_5160_1_108___stage___block_26_v_y)^(_q___pip_5160_1_108___stage___block_26_v_z);

_t___stage___block_2162_vnum0 = {_q___pip_5160_1_108___stage___block_26_v_z[0+:2],_q___pip_5160_1_108___stage___block_26_v_y[0+:2],_q___pip_5160_1_108___stage___block_26_v_x[0+:2]};

_t___stage___block_2162_vnum1 = {_q___pip_5160_1_108___stage___block_26_v_z[2+:2],_q___pip_5160_1_108___stage___block_26_v_y[2+:2],_q___pip_5160_1_108___stage___block_26_v_x[2+:2]};

_t___stage___block_2162_vnum2 = {_q___pip_5160_1_108___stage___block_26_v_z[4+:2],_q___pip_5160_1_108___stage___block_26_v_y[4+:2],_q___pip_5160_1_108___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_108___stage___block_6_inside&_w_tile[_t___stage___block_2162_vnum0+:1]&_w_tile[_t___stage___block_2162_vnum1+:1]&_w_tile[_t___stage___block_2162_vnum2+:1]) begin
// __block_2163
// __block_2165
_d___pip_5160_1_108___stage___block_6_clr = _t___stage___block_2162_tex;

_d___pip_5160_1_108___stage___block_6_dist = 188;

_d___pip_5160_1_108___stage___block_6_inside = 1;

// __block_2166
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2164
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2167
_t___block_2167_cmp_yx = _q___pip_5160_1_108___block_34_tm_y-_q___pip_5160_1_108___block_34_tm_x;

_t___block_2167_cmp_zx = _q___pip_5160_1_108___block_34_tm_z-_q___pip_5160_1_108___block_34_tm_x;

_t___block_2167_cmp_zy = _q___pip_5160_1_108___block_34_tm_z-_q___pip_5160_1_108___block_34_tm_y;

_t___block_2167_x_sel = ~_t___block_2167_cmp_yx[20+:1]&&~_t___block_2167_cmp_zx[20+:1];

_t___block_2167_y_sel = _t___block_2167_cmp_yx[20+:1]&&~_t___block_2167_cmp_zy[20+:1];

_t___block_2167_z_sel = _t___block_2167_cmp_zx[20+:1]&&_t___block_2167_cmp_zy[20+:1];

if (_t___block_2167_x_sel) begin
// __block_2168
// __block_2170
_d___pip_5160_1_108___stage___block_26_v_x = _q___pip_5160_1_108___stage___block_26_v_x+_q___pip_5160_1_108___stage___block_26_s_x;

_d___pip_5160_1_108___block_34_tm_x = _q___pip_5160_1_108___block_34_tm_x+_q___pip_5160_1_108___block_40_dt_x;

// __block_2171
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2169
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2172
if (_t___block_2167_y_sel) begin
// __block_2173
// __block_2175
_d___pip_5160_1_108___stage___block_26_v_y = _q___pip_5160_1_108___stage___block_26_v_y+_q___pip_5160_1_108___stage___block_26_s_y;

_d___pip_5160_1_108___block_34_tm_y = _q___pip_5160_1_108___block_34_tm_y+_q___pip_5160_1_108___block_40_dt_y;

// __block_2176
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2174
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2177
if (_t___block_2167_z_sel) begin
// __block_2178
// __block_2180
_d___pip_5160_1_108___stage___block_26_v_z = _q___pip_5160_1_108___stage___block_26_v_z+_q___pip_5160_1_108___stage___block_26_s_z;

_d___pip_5160_1_108___block_34_tm_z = _q___pip_5160_1_108___block_34_tm_z+_q___pip_5160_1_108___block_40_dt_z;

// __block_2181
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2179
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2182
// end of pipeline stage
_d__full_fsm___pip_5160_1_108 = 1;
_d__idx_fsm___pip_5160_1_108 = _t__stall_fsm___pip_5160_1_108 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_108 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 109
(* full_case *)
case (_q__idx_fsm___pip_5160_1_109)
1: begin
// __stage___block_2183
_t___stage___block_2183_tex = (_q___pip_5160_1_109___stage___block_26_v_x)^(_q___pip_5160_1_109___stage___block_26_v_y)^(_q___pip_5160_1_109___stage___block_26_v_z);

_t___stage___block_2183_vnum0 = {_q___pip_5160_1_109___stage___block_26_v_z[0+:2],_q___pip_5160_1_109___stage___block_26_v_y[0+:2],_q___pip_5160_1_109___stage___block_26_v_x[0+:2]};

_t___stage___block_2183_vnum1 = {_q___pip_5160_1_109___stage___block_26_v_z[2+:2],_q___pip_5160_1_109___stage___block_26_v_y[2+:2],_q___pip_5160_1_109___stage___block_26_v_x[2+:2]};

_t___stage___block_2183_vnum2 = {_q___pip_5160_1_109___stage___block_26_v_z[4+:2],_q___pip_5160_1_109___stage___block_26_v_y[4+:2],_q___pip_5160_1_109___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_109___stage___block_6_inside&_w_tile[_t___stage___block_2183_vnum0+:1]&_w_tile[_t___stage___block_2183_vnum1+:1]&_w_tile[_t___stage___block_2183_vnum2+:1]) begin
// __block_2184
// __block_2186
_d___pip_5160_1_109___stage___block_6_clr = _t___stage___block_2183_tex;

_d___pip_5160_1_109___stage___block_6_dist = 190;

_d___pip_5160_1_109___stage___block_6_inside = 1;

// __block_2187
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2185
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2188
_t___block_2188_cmp_yx = _q___pip_5160_1_109___block_34_tm_y-_q___pip_5160_1_109___block_34_tm_x;

_t___block_2188_cmp_zx = _q___pip_5160_1_109___block_34_tm_z-_q___pip_5160_1_109___block_34_tm_x;

_t___block_2188_cmp_zy = _q___pip_5160_1_109___block_34_tm_z-_q___pip_5160_1_109___block_34_tm_y;

_t___block_2188_x_sel = ~_t___block_2188_cmp_yx[20+:1]&&~_t___block_2188_cmp_zx[20+:1];

_t___block_2188_y_sel = _t___block_2188_cmp_yx[20+:1]&&~_t___block_2188_cmp_zy[20+:1];

_t___block_2188_z_sel = _t___block_2188_cmp_zx[20+:1]&&_t___block_2188_cmp_zy[20+:1];

if (_t___block_2188_x_sel) begin
// __block_2189
// __block_2191
_d___pip_5160_1_109___stage___block_26_v_x = _q___pip_5160_1_109___stage___block_26_v_x+_q___pip_5160_1_109___stage___block_26_s_x;

_d___pip_5160_1_109___block_34_tm_x = _q___pip_5160_1_109___block_34_tm_x+_q___pip_5160_1_109___block_40_dt_x;

// __block_2192
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2190
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2193
if (_t___block_2188_y_sel) begin
// __block_2194
// __block_2196
_d___pip_5160_1_109___stage___block_26_v_y = _q___pip_5160_1_109___stage___block_26_v_y+_q___pip_5160_1_109___stage___block_26_s_y;

_d___pip_5160_1_109___block_34_tm_y = _q___pip_5160_1_109___block_34_tm_y+_q___pip_5160_1_109___block_40_dt_y;

// __block_2197
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2195
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2198
if (_t___block_2188_z_sel) begin
// __block_2199
// __block_2201
_d___pip_5160_1_109___stage___block_26_v_z = _q___pip_5160_1_109___stage___block_26_v_z+_q___pip_5160_1_109___stage___block_26_s_z;

_d___pip_5160_1_109___block_34_tm_z = _q___pip_5160_1_109___block_34_tm_z+_q___pip_5160_1_109___block_40_dt_z;

// __block_2202
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2200
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2203
// end of pipeline stage
_d__full_fsm___pip_5160_1_109 = 1;
_d__idx_fsm___pip_5160_1_109 = _t__stall_fsm___pip_5160_1_109 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_109 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 110
(* full_case *)
case (_q__idx_fsm___pip_5160_1_110)
1: begin
// __stage___block_2204
_t___stage___block_2204_tex = (_q___pip_5160_1_110___stage___block_26_v_x)^(_q___pip_5160_1_110___stage___block_26_v_y)^(_q___pip_5160_1_110___stage___block_26_v_z);

_t___stage___block_2204_vnum0 = {_q___pip_5160_1_110___stage___block_26_v_z[0+:2],_q___pip_5160_1_110___stage___block_26_v_y[0+:2],_q___pip_5160_1_110___stage___block_26_v_x[0+:2]};

_t___stage___block_2204_vnum1 = {_q___pip_5160_1_110___stage___block_26_v_z[2+:2],_q___pip_5160_1_110___stage___block_26_v_y[2+:2],_q___pip_5160_1_110___stage___block_26_v_x[2+:2]};

_t___stage___block_2204_vnum2 = {_q___pip_5160_1_110___stage___block_26_v_z[4+:2],_q___pip_5160_1_110___stage___block_26_v_y[4+:2],_q___pip_5160_1_110___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_110___stage___block_6_inside&_w_tile[_t___stage___block_2204_vnum0+:1]&_w_tile[_t___stage___block_2204_vnum1+:1]&_w_tile[_t___stage___block_2204_vnum2+:1]) begin
// __block_2205
// __block_2207
_d___pip_5160_1_110___stage___block_6_clr = _t___stage___block_2204_tex;

_d___pip_5160_1_110___stage___block_6_dist = 192;

_d___pip_5160_1_110___stage___block_6_inside = 1;

// __block_2208
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2206
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2209
_t___block_2209_cmp_yx = _q___pip_5160_1_110___block_34_tm_y-_q___pip_5160_1_110___block_34_tm_x;

_t___block_2209_cmp_zx = _q___pip_5160_1_110___block_34_tm_z-_q___pip_5160_1_110___block_34_tm_x;

_t___block_2209_cmp_zy = _q___pip_5160_1_110___block_34_tm_z-_q___pip_5160_1_110___block_34_tm_y;

_t___block_2209_x_sel = ~_t___block_2209_cmp_yx[20+:1]&&~_t___block_2209_cmp_zx[20+:1];

_t___block_2209_y_sel = _t___block_2209_cmp_yx[20+:1]&&~_t___block_2209_cmp_zy[20+:1];

_t___block_2209_z_sel = _t___block_2209_cmp_zx[20+:1]&&_t___block_2209_cmp_zy[20+:1];

if (_t___block_2209_x_sel) begin
// __block_2210
// __block_2212
_d___pip_5160_1_110___stage___block_26_v_x = _q___pip_5160_1_110___stage___block_26_v_x+_q___pip_5160_1_110___stage___block_26_s_x;

_d___pip_5160_1_110___block_34_tm_x = _q___pip_5160_1_110___block_34_tm_x+_q___pip_5160_1_110___block_40_dt_x;

// __block_2213
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2211
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2214
if (_t___block_2209_y_sel) begin
// __block_2215
// __block_2217
_d___pip_5160_1_110___stage___block_26_v_y = _q___pip_5160_1_110___stage___block_26_v_y+_q___pip_5160_1_110___stage___block_26_s_y;

_d___pip_5160_1_110___block_34_tm_y = _q___pip_5160_1_110___block_34_tm_y+_q___pip_5160_1_110___block_40_dt_y;

// __block_2218
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2216
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2219
if (_t___block_2209_z_sel) begin
// __block_2220
// __block_2222
_d___pip_5160_1_110___stage___block_26_v_z = _q___pip_5160_1_110___stage___block_26_v_z+_q___pip_5160_1_110___stage___block_26_s_z;

_d___pip_5160_1_110___block_34_tm_z = _q___pip_5160_1_110___block_34_tm_z+_q___pip_5160_1_110___block_40_dt_z;

// __block_2223
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2221
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2224
// end of pipeline stage
_d__full_fsm___pip_5160_1_110 = 1;
_d__idx_fsm___pip_5160_1_110 = _t__stall_fsm___pip_5160_1_110 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_110 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 111
(* full_case *)
case (_q__idx_fsm___pip_5160_1_111)
1: begin
// __stage___block_2225
_t___stage___block_2225_tex = (_q___pip_5160_1_111___stage___block_26_v_x)^(_q___pip_5160_1_111___stage___block_26_v_y)^(_q___pip_5160_1_111___stage___block_26_v_z);

_t___stage___block_2225_vnum0 = {_q___pip_5160_1_111___stage___block_26_v_z[0+:2],_q___pip_5160_1_111___stage___block_26_v_y[0+:2],_q___pip_5160_1_111___stage___block_26_v_x[0+:2]};

_t___stage___block_2225_vnum1 = {_q___pip_5160_1_111___stage___block_26_v_z[2+:2],_q___pip_5160_1_111___stage___block_26_v_y[2+:2],_q___pip_5160_1_111___stage___block_26_v_x[2+:2]};

_t___stage___block_2225_vnum2 = {_q___pip_5160_1_111___stage___block_26_v_z[4+:2],_q___pip_5160_1_111___stage___block_26_v_y[4+:2],_q___pip_5160_1_111___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_111___stage___block_6_inside&_w_tile[_t___stage___block_2225_vnum0+:1]&_w_tile[_t___stage___block_2225_vnum1+:1]&_w_tile[_t___stage___block_2225_vnum2+:1]) begin
// __block_2226
// __block_2228
_d___pip_5160_1_111___stage___block_6_clr = _t___stage___block_2225_tex;

_d___pip_5160_1_111___stage___block_6_dist = 194;

_d___pip_5160_1_111___stage___block_6_inside = 1;

// __block_2229
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2227
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2230
_t___block_2230_cmp_yx = _q___pip_5160_1_111___block_34_tm_y-_q___pip_5160_1_111___block_34_tm_x;

_t___block_2230_cmp_zx = _q___pip_5160_1_111___block_34_tm_z-_q___pip_5160_1_111___block_34_tm_x;

_t___block_2230_cmp_zy = _q___pip_5160_1_111___block_34_tm_z-_q___pip_5160_1_111___block_34_tm_y;

_t___block_2230_x_sel = ~_t___block_2230_cmp_yx[20+:1]&&~_t___block_2230_cmp_zx[20+:1];

_t___block_2230_y_sel = _t___block_2230_cmp_yx[20+:1]&&~_t___block_2230_cmp_zy[20+:1];

_t___block_2230_z_sel = _t___block_2230_cmp_zx[20+:1]&&_t___block_2230_cmp_zy[20+:1];

if (_t___block_2230_x_sel) begin
// __block_2231
// __block_2233
_d___pip_5160_1_111___stage___block_26_v_x = _q___pip_5160_1_111___stage___block_26_v_x+_q___pip_5160_1_111___stage___block_26_s_x;

_d___pip_5160_1_111___block_34_tm_x = _q___pip_5160_1_111___block_34_tm_x+_q___pip_5160_1_111___block_40_dt_x;

// __block_2234
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2232
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2235
if (_t___block_2230_y_sel) begin
// __block_2236
// __block_2238
_d___pip_5160_1_111___stage___block_26_v_y = _q___pip_5160_1_111___stage___block_26_v_y+_q___pip_5160_1_111___stage___block_26_s_y;

_d___pip_5160_1_111___block_34_tm_y = _q___pip_5160_1_111___block_34_tm_y+_q___pip_5160_1_111___block_40_dt_y;

// __block_2239
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2237
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2240
if (_t___block_2230_z_sel) begin
// __block_2241
// __block_2243
_d___pip_5160_1_111___stage___block_26_v_z = _q___pip_5160_1_111___stage___block_26_v_z+_q___pip_5160_1_111___stage___block_26_s_z;

_d___pip_5160_1_111___block_34_tm_z = _q___pip_5160_1_111___block_34_tm_z+_q___pip_5160_1_111___block_40_dt_z;

// __block_2244
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2242
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2245
// end of pipeline stage
_d__full_fsm___pip_5160_1_111 = 1;
_d__idx_fsm___pip_5160_1_111 = _t__stall_fsm___pip_5160_1_111 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_111 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 112
(* full_case *)
case (_q__idx_fsm___pip_5160_1_112)
1: begin
// __stage___block_2246
_t___stage___block_2246_tex = (_q___pip_5160_1_112___stage___block_26_v_x)^(_q___pip_5160_1_112___stage___block_26_v_y)^(_q___pip_5160_1_112___stage___block_26_v_z);

_t___stage___block_2246_vnum0 = {_q___pip_5160_1_112___stage___block_26_v_z[0+:2],_q___pip_5160_1_112___stage___block_26_v_y[0+:2],_q___pip_5160_1_112___stage___block_26_v_x[0+:2]};

_t___stage___block_2246_vnum1 = {_q___pip_5160_1_112___stage___block_26_v_z[2+:2],_q___pip_5160_1_112___stage___block_26_v_y[2+:2],_q___pip_5160_1_112___stage___block_26_v_x[2+:2]};

_t___stage___block_2246_vnum2 = {_q___pip_5160_1_112___stage___block_26_v_z[4+:2],_q___pip_5160_1_112___stage___block_26_v_y[4+:2],_q___pip_5160_1_112___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_112___stage___block_6_inside&_w_tile[_t___stage___block_2246_vnum0+:1]&_w_tile[_t___stage___block_2246_vnum1+:1]&_w_tile[_t___stage___block_2246_vnum2+:1]) begin
// __block_2247
// __block_2249
_d___pip_5160_1_112___stage___block_6_clr = _t___stage___block_2246_tex;

_d___pip_5160_1_112___stage___block_6_dist = 196;

_d___pip_5160_1_112___stage___block_6_inside = 1;

// __block_2250
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2248
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2251
_t___block_2251_cmp_yx = _q___pip_5160_1_112___block_34_tm_y-_q___pip_5160_1_112___block_34_tm_x;

_t___block_2251_cmp_zx = _q___pip_5160_1_112___block_34_tm_z-_q___pip_5160_1_112___block_34_tm_x;

_t___block_2251_cmp_zy = _q___pip_5160_1_112___block_34_tm_z-_q___pip_5160_1_112___block_34_tm_y;

_t___block_2251_x_sel = ~_t___block_2251_cmp_yx[20+:1]&&~_t___block_2251_cmp_zx[20+:1];

_t___block_2251_y_sel = _t___block_2251_cmp_yx[20+:1]&&~_t___block_2251_cmp_zy[20+:1];

_t___block_2251_z_sel = _t___block_2251_cmp_zx[20+:1]&&_t___block_2251_cmp_zy[20+:1];

if (_t___block_2251_x_sel) begin
// __block_2252
// __block_2254
_d___pip_5160_1_112___stage___block_26_v_x = _q___pip_5160_1_112___stage___block_26_v_x+_q___pip_5160_1_112___stage___block_26_s_x;

_d___pip_5160_1_112___block_34_tm_x = _q___pip_5160_1_112___block_34_tm_x+_q___pip_5160_1_112___block_40_dt_x;

// __block_2255
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2253
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2256
if (_t___block_2251_y_sel) begin
// __block_2257
// __block_2259
_d___pip_5160_1_112___stage___block_26_v_y = _q___pip_5160_1_112___stage___block_26_v_y+_q___pip_5160_1_112___stage___block_26_s_y;

_d___pip_5160_1_112___block_34_tm_y = _q___pip_5160_1_112___block_34_tm_y+_q___pip_5160_1_112___block_40_dt_y;

// __block_2260
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2258
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2261
if (_t___block_2251_z_sel) begin
// __block_2262
// __block_2264
_d___pip_5160_1_112___stage___block_26_v_z = _q___pip_5160_1_112___stage___block_26_v_z+_q___pip_5160_1_112___stage___block_26_s_z;

_d___pip_5160_1_112___block_34_tm_z = _q___pip_5160_1_112___block_34_tm_z+_q___pip_5160_1_112___block_40_dt_z;

// __block_2265
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2263
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2266
// end of pipeline stage
_d__full_fsm___pip_5160_1_112 = 1;
_d__idx_fsm___pip_5160_1_112 = _t__stall_fsm___pip_5160_1_112 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_112 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 113
(* full_case *)
case (_q__idx_fsm___pip_5160_1_113)
1: begin
// __stage___block_2267
_t___stage___block_2267_tex = (_q___pip_5160_1_113___stage___block_26_v_x)^(_q___pip_5160_1_113___stage___block_26_v_y)^(_q___pip_5160_1_113___stage___block_26_v_z);

_t___stage___block_2267_vnum0 = {_q___pip_5160_1_113___stage___block_26_v_z[0+:2],_q___pip_5160_1_113___stage___block_26_v_y[0+:2],_q___pip_5160_1_113___stage___block_26_v_x[0+:2]};

_t___stage___block_2267_vnum1 = {_q___pip_5160_1_113___stage___block_26_v_z[2+:2],_q___pip_5160_1_113___stage___block_26_v_y[2+:2],_q___pip_5160_1_113___stage___block_26_v_x[2+:2]};

_t___stage___block_2267_vnum2 = {_q___pip_5160_1_113___stage___block_26_v_z[4+:2],_q___pip_5160_1_113___stage___block_26_v_y[4+:2],_q___pip_5160_1_113___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_113___stage___block_6_inside&_w_tile[_t___stage___block_2267_vnum0+:1]&_w_tile[_t___stage___block_2267_vnum1+:1]&_w_tile[_t___stage___block_2267_vnum2+:1]) begin
// __block_2268
// __block_2270
_d___pip_5160_1_113___stage___block_6_clr = _t___stage___block_2267_tex;

_d___pip_5160_1_113___stage___block_6_dist = 197;

_d___pip_5160_1_113___stage___block_6_inside = 1;

// __block_2271
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2269
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2272
_t___block_2272_cmp_yx = _q___pip_5160_1_113___block_34_tm_y-_q___pip_5160_1_113___block_34_tm_x;

_t___block_2272_cmp_zx = _q___pip_5160_1_113___block_34_tm_z-_q___pip_5160_1_113___block_34_tm_x;

_t___block_2272_cmp_zy = _q___pip_5160_1_113___block_34_tm_z-_q___pip_5160_1_113___block_34_tm_y;

_t___block_2272_x_sel = ~_t___block_2272_cmp_yx[20+:1]&&~_t___block_2272_cmp_zx[20+:1];

_t___block_2272_y_sel = _t___block_2272_cmp_yx[20+:1]&&~_t___block_2272_cmp_zy[20+:1];

_t___block_2272_z_sel = _t___block_2272_cmp_zx[20+:1]&&_t___block_2272_cmp_zy[20+:1];

if (_t___block_2272_x_sel) begin
// __block_2273
// __block_2275
_d___pip_5160_1_113___stage___block_26_v_x = _q___pip_5160_1_113___stage___block_26_v_x+_q___pip_5160_1_113___stage___block_26_s_x;

_d___pip_5160_1_113___block_34_tm_x = _q___pip_5160_1_113___block_34_tm_x+_q___pip_5160_1_113___block_40_dt_x;

// __block_2276
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2274
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2277
if (_t___block_2272_y_sel) begin
// __block_2278
// __block_2280
_d___pip_5160_1_113___stage___block_26_v_y = _q___pip_5160_1_113___stage___block_26_v_y+_q___pip_5160_1_113___stage___block_26_s_y;

_d___pip_5160_1_113___block_34_tm_y = _q___pip_5160_1_113___block_34_tm_y+_q___pip_5160_1_113___block_40_dt_y;

// __block_2281
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2279
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2282
if (_t___block_2272_z_sel) begin
// __block_2283
// __block_2285
_d___pip_5160_1_113___stage___block_26_v_z = _q___pip_5160_1_113___stage___block_26_v_z+_q___pip_5160_1_113___stage___block_26_s_z;

_d___pip_5160_1_113___block_34_tm_z = _q___pip_5160_1_113___block_34_tm_z+_q___pip_5160_1_113___block_40_dt_z;

// __block_2286
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2284
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2287
// end of pipeline stage
_d__full_fsm___pip_5160_1_113 = 1;
_d__idx_fsm___pip_5160_1_113 = _t__stall_fsm___pip_5160_1_113 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_113 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 114
(* full_case *)
case (_q__idx_fsm___pip_5160_1_114)
1: begin
// __stage___block_2288
_t___stage___block_2288_tex = (_q___pip_5160_1_114___stage___block_26_v_x)^(_q___pip_5160_1_114___stage___block_26_v_y)^(_q___pip_5160_1_114___stage___block_26_v_z);

_t___stage___block_2288_vnum0 = {_q___pip_5160_1_114___stage___block_26_v_z[0+:2],_q___pip_5160_1_114___stage___block_26_v_y[0+:2],_q___pip_5160_1_114___stage___block_26_v_x[0+:2]};

_t___stage___block_2288_vnum1 = {_q___pip_5160_1_114___stage___block_26_v_z[2+:2],_q___pip_5160_1_114___stage___block_26_v_y[2+:2],_q___pip_5160_1_114___stage___block_26_v_x[2+:2]};

_t___stage___block_2288_vnum2 = {_q___pip_5160_1_114___stage___block_26_v_z[4+:2],_q___pip_5160_1_114___stage___block_26_v_y[4+:2],_q___pip_5160_1_114___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_114___stage___block_6_inside&_w_tile[_t___stage___block_2288_vnum0+:1]&_w_tile[_t___stage___block_2288_vnum1+:1]&_w_tile[_t___stage___block_2288_vnum2+:1]) begin
// __block_2289
// __block_2291
_d___pip_5160_1_114___stage___block_6_clr = _t___stage___block_2288_tex;

_d___pip_5160_1_114___stage___block_6_dist = 199;

_d___pip_5160_1_114___stage___block_6_inside = 1;

// __block_2292
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2290
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2293
_t___block_2293_cmp_yx = _q___pip_5160_1_114___block_34_tm_y-_q___pip_5160_1_114___block_34_tm_x;

_t___block_2293_cmp_zx = _q___pip_5160_1_114___block_34_tm_z-_q___pip_5160_1_114___block_34_tm_x;

_t___block_2293_cmp_zy = _q___pip_5160_1_114___block_34_tm_z-_q___pip_5160_1_114___block_34_tm_y;

_t___block_2293_x_sel = ~_t___block_2293_cmp_yx[20+:1]&&~_t___block_2293_cmp_zx[20+:1];

_t___block_2293_y_sel = _t___block_2293_cmp_yx[20+:1]&&~_t___block_2293_cmp_zy[20+:1];

_t___block_2293_z_sel = _t___block_2293_cmp_zx[20+:1]&&_t___block_2293_cmp_zy[20+:1];

if (_t___block_2293_x_sel) begin
// __block_2294
// __block_2296
_d___pip_5160_1_114___stage___block_26_v_x = _q___pip_5160_1_114___stage___block_26_v_x+_q___pip_5160_1_114___stage___block_26_s_x;

_d___pip_5160_1_114___block_34_tm_x = _q___pip_5160_1_114___block_34_tm_x+_q___pip_5160_1_114___block_40_dt_x;

// __block_2297
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2295
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2298
if (_t___block_2293_y_sel) begin
// __block_2299
// __block_2301
_d___pip_5160_1_114___stage___block_26_v_y = _q___pip_5160_1_114___stage___block_26_v_y+_q___pip_5160_1_114___stage___block_26_s_y;

_d___pip_5160_1_114___block_34_tm_y = _q___pip_5160_1_114___block_34_tm_y+_q___pip_5160_1_114___block_40_dt_y;

// __block_2302
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2300
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2303
if (_t___block_2293_z_sel) begin
// __block_2304
// __block_2306
_d___pip_5160_1_114___stage___block_26_v_z = _q___pip_5160_1_114___stage___block_26_v_z+_q___pip_5160_1_114___stage___block_26_s_z;

_d___pip_5160_1_114___block_34_tm_z = _q___pip_5160_1_114___block_34_tm_z+_q___pip_5160_1_114___block_40_dt_z;

// __block_2307
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2305
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2308
// end of pipeline stage
_d__full_fsm___pip_5160_1_114 = 1;
_d__idx_fsm___pip_5160_1_114 = _t__stall_fsm___pip_5160_1_114 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_114 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 115
(* full_case *)
case (_q__idx_fsm___pip_5160_1_115)
1: begin
// __stage___block_2309
_t___stage___block_2309_tex = (_q___pip_5160_1_115___stage___block_26_v_x)^(_q___pip_5160_1_115___stage___block_26_v_y)^(_q___pip_5160_1_115___stage___block_26_v_z);

_t___stage___block_2309_vnum0 = {_q___pip_5160_1_115___stage___block_26_v_z[0+:2],_q___pip_5160_1_115___stage___block_26_v_y[0+:2],_q___pip_5160_1_115___stage___block_26_v_x[0+:2]};

_t___stage___block_2309_vnum1 = {_q___pip_5160_1_115___stage___block_26_v_z[2+:2],_q___pip_5160_1_115___stage___block_26_v_y[2+:2],_q___pip_5160_1_115___stage___block_26_v_x[2+:2]};

_t___stage___block_2309_vnum2 = {_q___pip_5160_1_115___stage___block_26_v_z[4+:2],_q___pip_5160_1_115___stage___block_26_v_y[4+:2],_q___pip_5160_1_115___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_115___stage___block_6_inside&_w_tile[_t___stage___block_2309_vnum0+:1]&_w_tile[_t___stage___block_2309_vnum1+:1]&_w_tile[_t___stage___block_2309_vnum2+:1]) begin
// __block_2310
// __block_2312
_d___pip_5160_1_115___stage___block_6_clr = _t___stage___block_2309_tex;

_d___pip_5160_1_115___stage___block_6_dist = 201;

_d___pip_5160_1_115___stage___block_6_inside = 1;

// __block_2313
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2311
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2314
_t___block_2314_cmp_yx = _q___pip_5160_1_115___block_34_tm_y-_q___pip_5160_1_115___block_34_tm_x;

_t___block_2314_cmp_zx = _q___pip_5160_1_115___block_34_tm_z-_q___pip_5160_1_115___block_34_tm_x;

_t___block_2314_cmp_zy = _q___pip_5160_1_115___block_34_tm_z-_q___pip_5160_1_115___block_34_tm_y;

_t___block_2314_x_sel = ~_t___block_2314_cmp_yx[20+:1]&&~_t___block_2314_cmp_zx[20+:1];

_t___block_2314_y_sel = _t___block_2314_cmp_yx[20+:1]&&~_t___block_2314_cmp_zy[20+:1];

_t___block_2314_z_sel = _t___block_2314_cmp_zx[20+:1]&&_t___block_2314_cmp_zy[20+:1];

if (_t___block_2314_x_sel) begin
// __block_2315
// __block_2317
_d___pip_5160_1_115___stage___block_26_v_x = _q___pip_5160_1_115___stage___block_26_v_x+_q___pip_5160_1_115___stage___block_26_s_x;

_d___pip_5160_1_115___block_34_tm_x = _q___pip_5160_1_115___block_34_tm_x+_q___pip_5160_1_115___block_40_dt_x;

// __block_2318
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2316
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2319
if (_t___block_2314_y_sel) begin
// __block_2320
// __block_2322
_d___pip_5160_1_115___stage___block_26_v_y = _q___pip_5160_1_115___stage___block_26_v_y+_q___pip_5160_1_115___stage___block_26_s_y;

_d___pip_5160_1_115___block_34_tm_y = _q___pip_5160_1_115___block_34_tm_y+_q___pip_5160_1_115___block_40_dt_y;

// __block_2323
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2321
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2324
if (_t___block_2314_z_sel) begin
// __block_2325
// __block_2327
_d___pip_5160_1_115___stage___block_26_v_z = _q___pip_5160_1_115___stage___block_26_v_z+_q___pip_5160_1_115___stage___block_26_s_z;

_d___pip_5160_1_115___block_34_tm_z = _q___pip_5160_1_115___block_34_tm_z+_q___pip_5160_1_115___block_40_dt_z;

// __block_2328
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2326
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2329
// end of pipeline stage
_d__full_fsm___pip_5160_1_115 = 1;
_d__idx_fsm___pip_5160_1_115 = _t__stall_fsm___pip_5160_1_115 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_115 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 116
(* full_case *)
case (_q__idx_fsm___pip_5160_1_116)
1: begin
// __stage___block_2330
_t___stage___block_2330_tex = (_q___pip_5160_1_116___stage___block_26_v_x)^(_q___pip_5160_1_116___stage___block_26_v_y)^(_q___pip_5160_1_116___stage___block_26_v_z);

_t___stage___block_2330_vnum0 = {_q___pip_5160_1_116___stage___block_26_v_z[0+:2],_q___pip_5160_1_116___stage___block_26_v_y[0+:2],_q___pip_5160_1_116___stage___block_26_v_x[0+:2]};

_t___stage___block_2330_vnum1 = {_q___pip_5160_1_116___stage___block_26_v_z[2+:2],_q___pip_5160_1_116___stage___block_26_v_y[2+:2],_q___pip_5160_1_116___stage___block_26_v_x[2+:2]};

_t___stage___block_2330_vnum2 = {_q___pip_5160_1_116___stage___block_26_v_z[4+:2],_q___pip_5160_1_116___stage___block_26_v_y[4+:2],_q___pip_5160_1_116___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_116___stage___block_6_inside&_w_tile[_t___stage___block_2330_vnum0+:1]&_w_tile[_t___stage___block_2330_vnum1+:1]&_w_tile[_t___stage___block_2330_vnum2+:1]) begin
// __block_2331
// __block_2333
_d___pip_5160_1_116___stage___block_6_clr = _t___stage___block_2330_tex;

_d___pip_5160_1_116___stage___block_6_dist = 203;

_d___pip_5160_1_116___stage___block_6_inside = 1;

// __block_2334
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2332
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2335
_t___block_2335_cmp_yx = _q___pip_5160_1_116___block_34_tm_y-_q___pip_5160_1_116___block_34_tm_x;

_t___block_2335_cmp_zx = _q___pip_5160_1_116___block_34_tm_z-_q___pip_5160_1_116___block_34_tm_x;

_t___block_2335_cmp_zy = _q___pip_5160_1_116___block_34_tm_z-_q___pip_5160_1_116___block_34_tm_y;

_t___block_2335_x_sel = ~_t___block_2335_cmp_yx[20+:1]&&~_t___block_2335_cmp_zx[20+:1];

_t___block_2335_y_sel = _t___block_2335_cmp_yx[20+:1]&&~_t___block_2335_cmp_zy[20+:1];

_t___block_2335_z_sel = _t___block_2335_cmp_zx[20+:1]&&_t___block_2335_cmp_zy[20+:1];

if (_t___block_2335_x_sel) begin
// __block_2336
// __block_2338
_d___pip_5160_1_116___stage___block_26_v_x = _q___pip_5160_1_116___stage___block_26_v_x+_q___pip_5160_1_116___stage___block_26_s_x;

_d___pip_5160_1_116___block_34_tm_x = _q___pip_5160_1_116___block_34_tm_x+_q___pip_5160_1_116___block_40_dt_x;

// __block_2339
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2337
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2340
if (_t___block_2335_y_sel) begin
// __block_2341
// __block_2343
_d___pip_5160_1_116___stage___block_26_v_y = _q___pip_5160_1_116___stage___block_26_v_y+_q___pip_5160_1_116___stage___block_26_s_y;

_d___pip_5160_1_116___block_34_tm_y = _q___pip_5160_1_116___block_34_tm_y+_q___pip_5160_1_116___block_40_dt_y;

// __block_2344
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2342
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2345
if (_t___block_2335_z_sel) begin
// __block_2346
// __block_2348
_d___pip_5160_1_116___stage___block_26_v_z = _q___pip_5160_1_116___stage___block_26_v_z+_q___pip_5160_1_116___stage___block_26_s_z;

_d___pip_5160_1_116___block_34_tm_z = _q___pip_5160_1_116___block_34_tm_z+_q___pip_5160_1_116___block_40_dt_z;

// __block_2349
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2347
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2350
// end of pipeline stage
_d__full_fsm___pip_5160_1_116 = 1;
_d__idx_fsm___pip_5160_1_116 = _t__stall_fsm___pip_5160_1_116 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_116 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 117
(* full_case *)
case (_q__idx_fsm___pip_5160_1_117)
1: begin
// __stage___block_2351
_t___stage___block_2351_tex = (_q___pip_5160_1_117___stage___block_26_v_x)^(_q___pip_5160_1_117___stage___block_26_v_y)^(_q___pip_5160_1_117___stage___block_26_v_z);

_t___stage___block_2351_vnum0 = {_q___pip_5160_1_117___stage___block_26_v_z[0+:2],_q___pip_5160_1_117___stage___block_26_v_y[0+:2],_q___pip_5160_1_117___stage___block_26_v_x[0+:2]};

_t___stage___block_2351_vnum1 = {_q___pip_5160_1_117___stage___block_26_v_z[2+:2],_q___pip_5160_1_117___stage___block_26_v_y[2+:2],_q___pip_5160_1_117___stage___block_26_v_x[2+:2]};

_t___stage___block_2351_vnum2 = {_q___pip_5160_1_117___stage___block_26_v_z[4+:2],_q___pip_5160_1_117___stage___block_26_v_y[4+:2],_q___pip_5160_1_117___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_117___stage___block_6_inside&_w_tile[_t___stage___block_2351_vnum0+:1]&_w_tile[_t___stage___block_2351_vnum1+:1]&_w_tile[_t___stage___block_2351_vnum2+:1]) begin
// __block_2352
// __block_2354
_d___pip_5160_1_117___stage___block_6_clr = _t___stage___block_2351_tex;

_d___pip_5160_1_117___stage___block_6_dist = 205;

_d___pip_5160_1_117___stage___block_6_inside = 1;

// __block_2355
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2353
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2356
_t___block_2356_cmp_yx = _q___pip_5160_1_117___block_34_tm_y-_q___pip_5160_1_117___block_34_tm_x;

_t___block_2356_cmp_zx = _q___pip_5160_1_117___block_34_tm_z-_q___pip_5160_1_117___block_34_tm_x;

_t___block_2356_cmp_zy = _q___pip_5160_1_117___block_34_tm_z-_q___pip_5160_1_117___block_34_tm_y;

_t___block_2356_x_sel = ~_t___block_2356_cmp_yx[20+:1]&&~_t___block_2356_cmp_zx[20+:1];

_t___block_2356_y_sel = _t___block_2356_cmp_yx[20+:1]&&~_t___block_2356_cmp_zy[20+:1];

_t___block_2356_z_sel = _t___block_2356_cmp_zx[20+:1]&&_t___block_2356_cmp_zy[20+:1];

if (_t___block_2356_x_sel) begin
// __block_2357
// __block_2359
_d___pip_5160_1_117___stage___block_26_v_x = _q___pip_5160_1_117___stage___block_26_v_x+_q___pip_5160_1_117___stage___block_26_s_x;

_d___pip_5160_1_117___block_34_tm_x = _q___pip_5160_1_117___block_34_tm_x+_q___pip_5160_1_117___block_40_dt_x;

// __block_2360
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2358
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2361
if (_t___block_2356_y_sel) begin
// __block_2362
// __block_2364
_d___pip_5160_1_117___stage___block_26_v_y = _q___pip_5160_1_117___stage___block_26_v_y+_q___pip_5160_1_117___stage___block_26_s_y;

_d___pip_5160_1_117___block_34_tm_y = _q___pip_5160_1_117___block_34_tm_y+_q___pip_5160_1_117___block_40_dt_y;

// __block_2365
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2363
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2366
if (_t___block_2356_z_sel) begin
// __block_2367
// __block_2369
_d___pip_5160_1_117___stage___block_26_v_z = _q___pip_5160_1_117___stage___block_26_v_z+_q___pip_5160_1_117___stage___block_26_s_z;

_d___pip_5160_1_117___block_34_tm_z = _q___pip_5160_1_117___block_34_tm_z+_q___pip_5160_1_117___block_40_dt_z;

// __block_2370
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2368
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2371
// end of pipeline stage
_d__full_fsm___pip_5160_1_117 = 1;
_d__idx_fsm___pip_5160_1_117 = _t__stall_fsm___pip_5160_1_117 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_117 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 118
(* full_case *)
case (_q__idx_fsm___pip_5160_1_118)
1: begin
// __stage___block_2372
_t___stage___block_2372_tex = (_q___pip_5160_1_118___stage___block_26_v_x)^(_q___pip_5160_1_118___stage___block_26_v_y)^(_q___pip_5160_1_118___stage___block_26_v_z);

_t___stage___block_2372_vnum0 = {_q___pip_5160_1_118___stage___block_26_v_z[0+:2],_q___pip_5160_1_118___stage___block_26_v_y[0+:2],_q___pip_5160_1_118___stage___block_26_v_x[0+:2]};

_t___stage___block_2372_vnum1 = {_q___pip_5160_1_118___stage___block_26_v_z[2+:2],_q___pip_5160_1_118___stage___block_26_v_y[2+:2],_q___pip_5160_1_118___stage___block_26_v_x[2+:2]};

_t___stage___block_2372_vnum2 = {_q___pip_5160_1_118___stage___block_26_v_z[4+:2],_q___pip_5160_1_118___stage___block_26_v_y[4+:2],_q___pip_5160_1_118___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_118___stage___block_6_inside&_w_tile[_t___stage___block_2372_vnum0+:1]&_w_tile[_t___stage___block_2372_vnum1+:1]&_w_tile[_t___stage___block_2372_vnum2+:1]) begin
// __block_2373
// __block_2375
_d___pip_5160_1_118___stage___block_6_clr = _t___stage___block_2372_tex;

_d___pip_5160_1_118___stage___block_6_dist = 207;

_d___pip_5160_1_118___stage___block_6_inside = 1;

// __block_2376
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2374
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2377
_t___block_2377_cmp_yx = _q___pip_5160_1_118___block_34_tm_y-_q___pip_5160_1_118___block_34_tm_x;

_t___block_2377_cmp_zx = _q___pip_5160_1_118___block_34_tm_z-_q___pip_5160_1_118___block_34_tm_x;

_t___block_2377_cmp_zy = _q___pip_5160_1_118___block_34_tm_z-_q___pip_5160_1_118___block_34_tm_y;

_t___block_2377_x_sel = ~_t___block_2377_cmp_yx[20+:1]&&~_t___block_2377_cmp_zx[20+:1];

_t___block_2377_y_sel = _t___block_2377_cmp_yx[20+:1]&&~_t___block_2377_cmp_zy[20+:1];

_t___block_2377_z_sel = _t___block_2377_cmp_zx[20+:1]&&_t___block_2377_cmp_zy[20+:1];

if (_t___block_2377_x_sel) begin
// __block_2378
// __block_2380
_d___pip_5160_1_118___stage___block_26_v_x = _q___pip_5160_1_118___stage___block_26_v_x+_q___pip_5160_1_118___stage___block_26_s_x;

_d___pip_5160_1_118___block_34_tm_x = _q___pip_5160_1_118___block_34_tm_x+_q___pip_5160_1_118___block_40_dt_x;

// __block_2381
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2379
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2382
if (_t___block_2377_y_sel) begin
// __block_2383
// __block_2385
_d___pip_5160_1_118___stage___block_26_v_y = _q___pip_5160_1_118___stage___block_26_v_y+_q___pip_5160_1_118___stage___block_26_s_y;

_d___pip_5160_1_118___block_34_tm_y = _q___pip_5160_1_118___block_34_tm_y+_q___pip_5160_1_118___block_40_dt_y;

// __block_2386
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2384
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2387
if (_t___block_2377_z_sel) begin
// __block_2388
// __block_2390
_d___pip_5160_1_118___stage___block_26_v_z = _q___pip_5160_1_118___stage___block_26_v_z+_q___pip_5160_1_118___stage___block_26_s_z;

_d___pip_5160_1_118___block_34_tm_z = _q___pip_5160_1_118___block_34_tm_z+_q___pip_5160_1_118___block_40_dt_z;

// __block_2391
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2389
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2392
// end of pipeline stage
_d__full_fsm___pip_5160_1_118 = 1;
_d__idx_fsm___pip_5160_1_118 = _t__stall_fsm___pip_5160_1_118 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_118 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 119
(* full_case *)
case (_q__idx_fsm___pip_5160_1_119)
1: begin
// __stage___block_2393
_t___stage___block_2393_tex = (_q___pip_5160_1_119___stage___block_26_v_x)^(_q___pip_5160_1_119___stage___block_26_v_y)^(_q___pip_5160_1_119___stage___block_26_v_z);

_t___stage___block_2393_vnum0 = {_q___pip_5160_1_119___stage___block_26_v_z[0+:2],_q___pip_5160_1_119___stage___block_26_v_y[0+:2],_q___pip_5160_1_119___stage___block_26_v_x[0+:2]};

_t___stage___block_2393_vnum1 = {_q___pip_5160_1_119___stage___block_26_v_z[2+:2],_q___pip_5160_1_119___stage___block_26_v_y[2+:2],_q___pip_5160_1_119___stage___block_26_v_x[2+:2]};

_t___stage___block_2393_vnum2 = {_q___pip_5160_1_119___stage___block_26_v_z[4+:2],_q___pip_5160_1_119___stage___block_26_v_y[4+:2],_q___pip_5160_1_119___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_119___stage___block_6_inside&_w_tile[_t___stage___block_2393_vnum0+:1]&_w_tile[_t___stage___block_2393_vnum1+:1]&_w_tile[_t___stage___block_2393_vnum2+:1]) begin
// __block_2394
// __block_2396
_d___pip_5160_1_119___stage___block_6_clr = _t___stage___block_2393_tex;

_d___pip_5160_1_119___stage___block_6_dist = 209;

_d___pip_5160_1_119___stage___block_6_inside = 1;

// __block_2397
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2395
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2398
_t___block_2398_cmp_yx = _q___pip_5160_1_119___block_34_tm_y-_q___pip_5160_1_119___block_34_tm_x;

_t___block_2398_cmp_zx = _q___pip_5160_1_119___block_34_tm_z-_q___pip_5160_1_119___block_34_tm_x;

_t___block_2398_cmp_zy = _q___pip_5160_1_119___block_34_tm_z-_q___pip_5160_1_119___block_34_tm_y;

_t___block_2398_x_sel = ~_t___block_2398_cmp_yx[20+:1]&&~_t___block_2398_cmp_zx[20+:1];

_t___block_2398_y_sel = _t___block_2398_cmp_yx[20+:1]&&~_t___block_2398_cmp_zy[20+:1];

_t___block_2398_z_sel = _t___block_2398_cmp_zx[20+:1]&&_t___block_2398_cmp_zy[20+:1];

if (_t___block_2398_x_sel) begin
// __block_2399
// __block_2401
_d___pip_5160_1_119___stage___block_26_v_x = _q___pip_5160_1_119___stage___block_26_v_x+_q___pip_5160_1_119___stage___block_26_s_x;

_d___pip_5160_1_119___block_34_tm_x = _q___pip_5160_1_119___block_34_tm_x+_q___pip_5160_1_119___block_40_dt_x;

// __block_2402
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2400
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2403
if (_t___block_2398_y_sel) begin
// __block_2404
// __block_2406
_d___pip_5160_1_119___stage___block_26_v_y = _q___pip_5160_1_119___stage___block_26_v_y+_q___pip_5160_1_119___stage___block_26_s_y;

_d___pip_5160_1_119___block_34_tm_y = _q___pip_5160_1_119___block_34_tm_y+_q___pip_5160_1_119___block_40_dt_y;

// __block_2407
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2405
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2408
if (_t___block_2398_z_sel) begin
// __block_2409
// __block_2411
_d___pip_5160_1_119___stage___block_26_v_z = _q___pip_5160_1_119___stage___block_26_v_z+_q___pip_5160_1_119___stage___block_26_s_z;

_d___pip_5160_1_119___block_34_tm_z = _q___pip_5160_1_119___block_34_tm_z+_q___pip_5160_1_119___block_40_dt_z;

// __block_2412
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2410
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2413
// end of pipeline stage
_d__full_fsm___pip_5160_1_119 = 1;
_d__idx_fsm___pip_5160_1_119 = _t__stall_fsm___pip_5160_1_119 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_119 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 120
(* full_case *)
case (_q__idx_fsm___pip_5160_1_120)
1: begin
// __stage___block_2414
_t___stage___block_2414_tex = (_q___pip_5160_1_120___stage___block_26_v_x)^(_q___pip_5160_1_120___stage___block_26_v_y)^(_q___pip_5160_1_120___stage___block_26_v_z);

_t___stage___block_2414_vnum0 = {_q___pip_5160_1_120___stage___block_26_v_z[0+:2],_q___pip_5160_1_120___stage___block_26_v_y[0+:2],_q___pip_5160_1_120___stage___block_26_v_x[0+:2]};

_t___stage___block_2414_vnum1 = {_q___pip_5160_1_120___stage___block_26_v_z[2+:2],_q___pip_5160_1_120___stage___block_26_v_y[2+:2],_q___pip_5160_1_120___stage___block_26_v_x[2+:2]};

_t___stage___block_2414_vnum2 = {_q___pip_5160_1_120___stage___block_26_v_z[4+:2],_q___pip_5160_1_120___stage___block_26_v_y[4+:2],_q___pip_5160_1_120___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_120___stage___block_6_inside&_w_tile[_t___stage___block_2414_vnum0+:1]&_w_tile[_t___stage___block_2414_vnum1+:1]&_w_tile[_t___stage___block_2414_vnum2+:1]) begin
// __block_2415
// __block_2417
_d___pip_5160_1_120___stage___block_6_clr = _t___stage___block_2414_tex;

_d___pip_5160_1_120___stage___block_6_dist = 210;

_d___pip_5160_1_120___stage___block_6_inside = 1;

// __block_2418
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2416
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2419
_t___block_2419_cmp_yx = _q___pip_5160_1_120___block_34_tm_y-_q___pip_5160_1_120___block_34_tm_x;

_t___block_2419_cmp_zx = _q___pip_5160_1_120___block_34_tm_z-_q___pip_5160_1_120___block_34_tm_x;

_t___block_2419_cmp_zy = _q___pip_5160_1_120___block_34_tm_z-_q___pip_5160_1_120___block_34_tm_y;

_t___block_2419_x_sel = ~_t___block_2419_cmp_yx[20+:1]&&~_t___block_2419_cmp_zx[20+:1];

_t___block_2419_y_sel = _t___block_2419_cmp_yx[20+:1]&&~_t___block_2419_cmp_zy[20+:1];

_t___block_2419_z_sel = _t___block_2419_cmp_zx[20+:1]&&_t___block_2419_cmp_zy[20+:1];

if (_t___block_2419_x_sel) begin
// __block_2420
// __block_2422
_d___pip_5160_1_120___stage___block_26_v_x = _q___pip_5160_1_120___stage___block_26_v_x+_q___pip_5160_1_120___stage___block_26_s_x;

_d___pip_5160_1_120___block_34_tm_x = _q___pip_5160_1_120___block_34_tm_x+_q___pip_5160_1_120___block_40_dt_x;

// __block_2423
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2421
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2424
if (_t___block_2419_y_sel) begin
// __block_2425
// __block_2427
_d___pip_5160_1_120___stage___block_26_v_y = _q___pip_5160_1_120___stage___block_26_v_y+_q___pip_5160_1_120___stage___block_26_s_y;

_d___pip_5160_1_120___block_34_tm_y = _q___pip_5160_1_120___block_34_tm_y+_q___pip_5160_1_120___block_40_dt_y;

// __block_2428
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2426
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2429
if (_t___block_2419_z_sel) begin
// __block_2430
// __block_2432
_d___pip_5160_1_120___stage___block_26_v_z = _q___pip_5160_1_120___stage___block_26_v_z+_q___pip_5160_1_120___stage___block_26_s_z;

_d___pip_5160_1_120___block_34_tm_z = _q___pip_5160_1_120___block_34_tm_z+_q___pip_5160_1_120___block_40_dt_z;

// __block_2433
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2431
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2434
// end of pipeline stage
_d__full_fsm___pip_5160_1_120 = 1;
_d__idx_fsm___pip_5160_1_120 = _t__stall_fsm___pip_5160_1_120 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_120 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 121
(* full_case *)
case (_q__idx_fsm___pip_5160_1_121)
1: begin
// __stage___block_2435
_t___stage___block_2435_tex = (_q___pip_5160_1_121___stage___block_26_v_x)^(_q___pip_5160_1_121___stage___block_26_v_y)^(_q___pip_5160_1_121___stage___block_26_v_z);

_t___stage___block_2435_vnum0 = {_q___pip_5160_1_121___stage___block_26_v_z[0+:2],_q___pip_5160_1_121___stage___block_26_v_y[0+:2],_q___pip_5160_1_121___stage___block_26_v_x[0+:2]};

_t___stage___block_2435_vnum1 = {_q___pip_5160_1_121___stage___block_26_v_z[2+:2],_q___pip_5160_1_121___stage___block_26_v_y[2+:2],_q___pip_5160_1_121___stage___block_26_v_x[2+:2]};

_t___stage___block_2435_vnum2 = {_q___pip_5160_1_121___stage___block_26_v_z[4+:2],_q___pip_5160_1_121___stage___block_26_v_y[4+:2],_q___pip_5160_1_121___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_121___stage___block_6_inside&_w_tile[_t___stage___block_2435_vnum0+:1]&_w_tile[_t___stage___block_2435_vnum1+:1]&_w_tile[_t___stage___block_2435_vnum2+:1]) begin
// __block_2436
// __block_2438
_d___pip_5160_1_121___stage___block_6_clr = _t___stage___block_2435_tex;

_d___pip_5160_1_121___stage___block_6_dist = 212;

_d___pip_5160_1_121___stage___block_6_inside = 1;

// __block_2439
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2437
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2440
_t___block_2440_cmp_yx = _q___pip_5160_1_121___block_34_tm_y-_q___pip_5160_1_121___block_34_tm_x;

_t___block_2440_cmp_zx = _q___pip_5160_1_121___block_34_tm_z-_q___pip_5160_1_121___block_34_tm_x;

_t___block_2440_cmp_zy = _q___pip_5160_1_121___block_34_tm_z-_q___pip_5160_1_121___block_34_tm_y;

_t___block_2440_x_sel = ~_t___block_2440_cmp_yx[20+:1]&&~_t___block_2440_cmp_zx[20+:1];

_t___block_2440_y_sel = _t___block_2440_cmp_yx[20+:1]&&~_t___block_2440_cmp_zy[20+:1];

_t___block_2440_z_sel = _t___block_2440_cmp_zx[20+:1]&&_t___block_2440_cmp_zy[20+:1];

if (_t___block_2440_x_sel) begin
// __block_2441
// __block_2443
_d___pip_5160_1_121___stage___block_26_v_x = _q___pip_5160_1_121___stage___block_26_v_x+_q___pip_5160_1_121___stage___block_26_s_x;

_d___pip_5160_1_121___block_34_tm_x = _q___pip_5160_1_121___block_34_tm_x+_q___pip_5160_1_121___block_40_dt_x;

// __block_2444
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2442
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2445
if (_t___block_2440_y_sel) begin
// __block_2446
// __block_2448
_d___pip_5160_1_121___stage___block_26_v_y = _q___pip_5160_1_121___stage___block_26_v_y+_q___pip_5160_1_121___stage___block_26_s_y;

_d___pip_5160_1_121___block_34_tm_y = _q___pip_5160_1_121___block_34_tm_y+_q___pip_5160_1_121___block_40_dt_y;

// __block_2449
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2447
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2450
if (_t___block_2440_z_sel) begin
// __block_2451
// __block_2453
_d___pip_5160_1_121___stage___block_26_v_z = _q___pip_5160_1_121___stage___block_26_v_z+_q___pip_5160_1_121___stage___block_26_s_z;

_d___pip_5160_1_121___block_34_tm_z = _q___pip_5160_1_121___block_34_tm_z+_q___pip_5160_1_121___block_40_dt_z;

// __block_2454
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2452
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2455
// end of pipeline stage
_d__full_fsm___pip_5160_1_121 = 1;
_d__idx_fsm___pip_5160_1_121 = _t__stall_fsm___pip_5160_1_121 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_121 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 122
(* full_case *)
case (_q__idx_fsm___pip_5160_1_122)
1: begin
// __stage___block_2456
_t___stage___block_2456_tex = (_q___pip_5160_1_122___stage___block_26_v_x)^(_q___pip_5160_1_122___stage___block_26_v_y)^(_q___pip_5160_1_122___stage___block_26_v_z);

_t___stage___block_2456_vnum0 = {_q___pip_5160_1_122___stage___block_26_v_z[0+:2],_q___pip_5160_1_122___stage___block_26_v_y[0+:2],_q___pip_5160_1_122___stage___block_26_v_x[0+:2]};

_t___stage___block_2456_vnum1 = {_q___pip_5160_1_122___stage___block_26_v_z[2+:2],_q___pip_5160_1_122___stage___block_26_v_y[2+:2],_q___pip_5160_1_122___stage___block_26_v_x[2+:2]};

_t___stage___block_2456_vnum2 = {_q___pip_5160_1_122___stage___block_26_v_z[4+:2],_q___pip_5160_1_122___stage___block_26_v_y[4+:2],_q___pip_5160_1_122___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_122___stage___block_6_inside&_w_tile[_t___stage___block_2456_vnum0+:1]&_w_tile[_t___stage___block_2456_vnum1+:1]&_w_tile[_t___stage___block_2456_vnum2+:1]) begin
// __block_2457
// __block_2459
_d___pip_5160_1_122___stage___block_6_clr = _t___stage___block_2456_tex;

_d___pip_5160_1_122___stage___block_6_dist = 214;

_d___pip_5160_1_122___stage___block_6_inside = 1;

// __block_2460
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2458
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2461
_t___block_2461_cmp_yx = _q___pip_5160_1_122___block_34_tm_y-_q___pip_5160_1_122___block_34_tm_x;

_t___block_2461_cmp_zx = _q___pip_5160_1_122___block_34_tm_z-_q___pip_5160_1_122___block_34_tm_x;

_t___block_2461_cmp_zy = _q___pip_5160_1_122___block_34_tm_z-_q___pip_5160_1_122___block_34_tm_y;

_t___block_2461_x_sel = ~_t___block_2461_cmp_yx[20+:1]&&~_t___block_2461_cmp_zx[20+:1];

_t___block_2461_y_sel = _t___block_2461_cmp_yx[20+:1]&&~_t___block_2461_cmp_zy[20+:1];

_t___block_2461_z_sel = _t___block_2461_cmp_zx[20+:1]&&_t___block_2461_cmp_zy[20+:1];

if (_t___block_2461_x_sel) begin
// __block_2462
// __block_2464
_d___pip_5160_1_122___stage___block_26_v_x = _q___pip_5160_1_122___stage___block_26_v_x+_q___pip_5160_1_122___stage___block_26_s_x;

_d___pip_5160_1_122___block_34_tm_x = _q___pip_5160_1_122___block_34_tm_x+_q___pip_5160_1_122___block_40_dt_x;

// __block_2465
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2463
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2466
if (_t___block_2461_y_sel) begin
// __block_2467
// __block_2469
_d___pip_5160_1_122___stage___block_26_v_y = _q___pip_5160_1_122___stage___block_26_v_y+_q___pip_5160_1_122___stage___block_26_s_y;

_d___pip_5160_1_122___block_34_tm_y = _q___pip_5160_1_122___block_34_tm_y+_q___pip_5160_1_122___block_40_dt_y;

// __block_2470
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2468
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2471
if (_t___block_2461_z_sel) begin
// __block_2472
// __block_2474
_d___pip_5160_1_122___stage___block_26_v_z = _q___pip_5160_1_122___stage___block_26_v_z+_q___pip_5160_1_122___stage___block_26_s_z;

_d___pip_5160_1_122___block_34_tm_z = _q___pip_5160_1_122___block_34_tm_z+_q___pip_5160_1_122___block_40_dt_z;

// __block_2475
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2473
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2476
// end of pipeline stage
_d__full_fsm___pip_5160_1_122 = 1;
_d__idx_fsm___pip_5160_1_122 = _t__stall_fsm___pip_5160_1_122 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_122 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 123
(* full_case *)
case (_q__idx_fsm___pip_5160_1_123)
1: begin
// __stage___block_2477
_t___stage___block_2477_tex = (_q___pip_5160_1_123___stage___block_26_v_x)^(_q___pip_5160_1_123___stage___block_26_v_y)^(_q___pip_5160_1_123___stage___block_26_v_z);

_t___stage___block_2477_vnum0 = {_q___pip_5160_1_123___stage___block_26_v_z[0+:2],_q___pip_5160_1_123___stage___block_26_v_y[0+:2],_q___pip_5160_1_123___stage___block_26_v_x[0+:2]};

_t___stage___block_2477_vnum1 = {_q___pip_5160_1_123___stage___block_26_v_z[2+:2],_q___pip_5160_1_123___stage___block_26_v_y[2+:2],_q___pip_5160_1_123___stage___block_26_v_x[2+:2]};

_t___stage___block_2477_vnum2 = {_q___pip_5160_1_123___stage___block_26_v_z[4+:2],_q___pip_5160_1_123___stage___block_26_v_y[4+:2],_q___pip_5160_1_123___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_123___stage___block_6_inside&_w_tile[_t___stage___block_2477_vnum0+:1]&_w_tile[_t___stage___block_2477_vnum1+:1]&_w_tile[_t___stage___block_2477_vnum2+:1]) begin
// __block_2478
// __block_2480
_d___pip_5160_1_123___stage___block_6_clr = _t___stage___block_2477_tex;

_d___pip_5160_1_123___stage___block_6_dist = 216;

_d___pip_5160_1_123___stage___block_6_inside = 1;

// __block_2481
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2479
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2482
_t___block_2482_cmp_yx = _q___pip_5160_1_123___block_34_tm_y-_q___pip_5160_1_123___block_34_tm_x;

_t___block_2482_cmp_zx = _q___pip_5160_1_123___block_34_tm_z-_q___pip_5160_1_123___block_34_tm_x;

_t___block_2482_cmp_zy = _q___pip_5160_1_123___block_34_tm_z-_q___pip_5160_1_123___block_34_tm_y;

_t___block_2482_x_sel = ~_t___block_2482_cmp_yx[20+:1]&&~_t___block_2482_cmp_zx[20+:1];

_t___block_2482_y_sel = _t___block_2482_cmp_yx[20+:1]&&~_t___block_2482_cmp_zy[20+:1];

_t___block_2482_z_sel = _t___block_2482_cmp_zx[20+:1]&&_t___block_2482_cmp_zy[20+:1];

if (_t___block_2482_x_sel) begin
// __block_2483
// __block_2485
_d___pip_5160_1_123___stage___block_26_v_x = _q___pip_5160_1_123___stage___block_26_v_x+_q___pip_5160_1_123___stage___block_26_s_x;

_d___pip_5160_1_123___block_34_tm_x = _q___pip_5160_1_123___block_34_tm_x+_q___pip_5160_1_123___block_40_dt_x;

// __block_2486
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2484
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2487
if (_t___block_2482_y_sel) begin
// __block_2488
// __block_2490
_d___pip_5160_1_123___stage___block_26_v_y = _q___pip_5160_1_123___stage___block_26_v_y+_q___pip_5160_1_123___stage___block_26_s_y;

_d___pip_5160_1_123___block_34_tm_y = _q___pip_5160_1_123___block_34_tm_y+_q___pip_5160_1_123___block_40_dt_y;

// __block_2491
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2489
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2492
if (_t___block_2482_z_sel) begin
// __block_2493
// __block_2495
_d___pip_5160_1_123___stage___block_26_v_z = _q___pip_5160_1_123___stage___block_26_v_z+_q___pip_5160_1_123___stage___block_26_s_z;

_d___pip_5160_1_123___block_34_tm_z = _q___pip_5160_1_123___block_34_tm_z+_q___pip_5160_1_123___block_40_dt_z;

// __block_2496
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2494
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2497
// end of pipeline stage
_d__full_fsm___pip_5160_1_123 = 1;
_d__idx_fsm___pip_5160_1_123 = _t__stall_fsm___pip_5160_1_123 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_123 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 124
(* full_case *)
case (_q__idx_fsm___pip_5160_1_124)
1: begin
// __stage___block_2498
_t___stage___block_2498_tex = (_q___pip_5160_1_124___stage___block_26_v_x)^(_q___pip_5160_1_124___stage___block_26_v_y)^(_q___pip_5160_1_124___stage___block_26_v_z);

_t___stage___block_2498_vnum0 = {_q___pip_5160_1_124___stage___block_26_v_z[0+:2],_q___pip_5160_1_124___stage___block_26_v_y[0+:2],_q___pip_5160_1_124___stage___block_26_v_x[0+:2]};

_t___stage___block_2498_vnum1 = {_q___pip_5160_1_124___stage___block_26_v_z[2+:2],_q___pip_5160_1_124___stage___block_26_v_y[2+:2],_q___pip_5160_1_124___stage___block_26_v_x[2+:2]};

_t___stage___block_2498_vnum2 = {_q___pip_5160_1_124___stage___block_26_v_z[4+:2],_q___pip_5160_1_124___stage___block_26_v_y[4+:2],_q___pip_5160_1_124___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_124___stage___block_6_inside&_w_tile[_t___stage___block_2498_vnum0+:1]&_w_tile[_t___stage___block_2498_vnum1+:1]&_w_tile[_t___stage___block_2498_vnum2+:1]) begin
// __block_2499
// __block_2501
_d___pip_5160_1_124___stage___block_6_clr = _t___stage___block_2498_tex;

_d___pip_5160_1_124___stage___block_6_dist = 218;

_d___pip_5160_1_124___stage___block_6_inside = 1;

// __block_2502
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2500
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2503
_t___block_2503_cmp_yx = _q___pip_5160_1_124___block_34_tm_y-_q___pip_5160_1_124___block_34_tm_x;

_t___block_2503_cmp_zx = _q___pip_5160_1_124___block_34_tm_z-_q___pip_5160_1_124___block_34_tm_x;

_t___block_2503_cmp_zy = _q___pip_5160_1_124___block_34_tm_z-_q___pip_5160_1_124___block_34_tm_y;

_t___block_2503_x_sel = ~_t___block_2503_cmp_yx[20+:1]&&~_t___block_2503_cmp_zx[20+:1];

_t___block_2503_y_sel = _t___block_2503_cmp_yx[20+:1]&&~_t___block_2503_cmp_zy[20+:1];

_t___block_2503_z_sel = _t___block_2503_cmp_zx[20+:1]&&_t___block_2503_cmp_zy[20+:1];

if (_t___block_2503_x_sel) begin
// __block_2504
// __block_2506
_d___pip_5160_1_124___stage___block_26_v_x = _q___pip_5160_1_124___stage___block_26_v_x+_q___pip_5160_1_124___stage___block_26_s_x;

_d___pip_5160_1_124___block_34_tm_x = _q___pip_5160_1_124___block_34_tm_x+_q___pip_5160_1_124___block_40_dt_x;

// __block_2507
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2505
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2508
if (_t___block_2503_y_sel) begin
// __block_2509
// __block_2511
_d___pip_5160_1_124___stage___block_26_v_y = _q___pip_5160_1_124___stage___block_26_v_y+_q___pip_5160_1_124___stage___block_26_s_y;

_d___pip_5160_1_124___block_34_tm_y = _q___pip_5160_1_124___block_34_tm_y+_q___pip_5160_1_124___block_40_dt_y;

// __block_2512
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2510
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2513
if (_t___block_2503_z_sel) begin
// __block_2514
// __block_2516
_d___pip_5160_1_124___stage___block_26_v_z = _q___pip_5160_1_124___stage___block_26_v_z+_q___pip_5160_1_124___stage___block_26_s_z;

_d___pip_5160_1_124___block_34_tm_z = _q___pip_5160_1_124___block_34_tm_z+_q___pip_5160_1_124___block_40_dt_z;

// __block_2517
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2515
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2518
// end of pipeline stage
_d__full_fsm___pip_5160_1_124 = 1;
_d__idx_fsm___pip_5160_1_124 = _t__stall_fsm___pip_5160_1_124 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_124 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 125
(* full_case *)
case (_q__idx_fsm___pip_5160_1_125)
1: begin
// __stage___block_2519
_t___stage___block_2519_tex = (_q___pip_5160_1_125___stage___block_26_v_x)^(_q___pip_5160_1_125___stage___block_26_v_y)^(_q___pip_5160_1_125___stage___block_26_v_z);

_t___stage___block_2519_vnum0 = {_q___pip_5160_1_125___stage___block_26_v_z[0+:2],_q___pip_5160_1_125___stage___block_26_v_y[0+:2],_q___pip_5160_1_125___stage___block_26_v_x[0+:2]};

_t___stage___block_2519_vnum1 = {_q___pip_5160_1_125___stage___block_26_v_z[2+:2],_q___pip_5160_1_125___stage___block_26_v_y[2+:2],_q___pip_5160_1_125___stage___block_26_v_x[2+:2]};

_t___stage___block_2519_vnum2 = {_q___pip_5160_1_125___stage___block_26_v_z[4+:2],_q___pip_5160_1_125___stage___block_26_v_y[4+:2],_q___pip_5160_1_125___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_125___stage___block_6_inside&_w_tile[_t___stage___block_2519_vnum0+:1]&_w_tile[_t___stage___block_2519_vnum1+:1]&_w_tile[_t___stage___block_2519_vnum2+:1]) begin
// __block_2520
// __block_2522
_d___pip_5160_1_125___stage___block_6_clr = _t___stage___block_2519_tex;

_d___pip_5160_1_125___stage___block_6_dist = 220;

_d___pip_5160_1_125___stage___block_6_inside = 1;

// __block_2523
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2521
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2524
_t___block_2524_cmp_yx = _q___pip_5160_1_125___block_34_tm_y-_q___pip_5160_1_125___block_34_tm_x;

_t___block_2524_cmp_zx = _q___pip_5160_1_125___block_34_tm_z-_q___pip_5160_1_125___block_34_tm_x;

_t___block_2524_cmp_zy = _q___pip_5160_1_125___block_34_tm_z-_q___pip_5160_1_125___block_34_tm_y;

_t___block_2524_x_sel = ~_t___block_2524_cmp_yx[20+:1]&&~_t___block_2524_cmp_zx[20+:1];

_t___block_2524_y_sel = _t___block_2524_cmp_yx[20+:1]&&~_t___block_2524_cmp_zy[20+:1];

_t___block_2524_z_sel = _t___block_2524_cmp_zx[20+:1]&&_t___block_2524_cmp_zy[20+:1];

if (_t___block_2524_x_sel) begin
// __block_2525
// __block_2527
_d___pip_5160_1_125___stage___block_26_v_x = _q___pip_5160_1_125___stage___block_26_v_x+_q___pip_5160_1_125___stage___block_26_s_x;

_d___pip_5160_1_125___block_34_tm_x = _q___pip_5160_1_125___block_34_tm_x+_q___pip_5160_1_125___block_40_dt_x;

// __block_2528
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2526
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2529
if (_t___block_2524_y_sel) begin
// __block_2530
// __block_2532
_d___pip_5160_1_125___stage___block_26_v_y = _q___pip_5160_1_125___stage___block_26_v_y+_q___pip_5160_1_125___stage___block_26_s_y;

_d___pip_5160_1_125___block_34_tm_y = _q___pip_5160_1_125___block_34_tm_y+_q___pip_5160_1_125___block_40_dt_y;

// __block_2533
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2531
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2534
if (_t___block_2524_z_sel) begin
// __block_2535
// __block_2537
_d___pip_5160_1_125___stage___block_26_v_z = _q___pip_5160_1_125___stage___block_26_v_z+_q___pip_5160_1_125___stage___block_26_s_z;

_d___pip_5160_1_125___block_34_tm_z = _q___pip_5160_1_125___block_34_tm_z+_q___pip_5160_1_125___block_40_dt_z;

// __block_2538
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2536
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2539
// end of pipeline stage
_d__full_fsm___pip_5160_1_125 = 1;
_d__idx_fsm___pip_5160_1_125 = _t__stall_fsm___pip_5160_1_125 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_125 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 126
(* full_case *)
case (_q__idx_fsm___pip_5160_1_126)
1: begin
// __stage___block_2540
_t___stage___block_2540_tex = (_q___pip_5160_1_126___stage___block_26_v_x)^(_q___pip_5160_1_126___stage___block_26_v_y)^(_q___pip_5160_1_126___stage___block_26_v_z);

_t___stage___block_2540_vnum0 = {_q___pip_5160_1_126___stage___block_26_v_z[0+:2],_q___pip_5160_1_126___stage___block_26_v_y[0+:2],_q___pip_5160_1_126___stage___block_26_v_x[0+:2]};

_t___stage___block_2540_vnum1 = {_q___pip_5160_1_126___stage___block_26_v_z[2+:2],_q___pip_5160_1_126___stage___block_26_v_y[2+:2],_q___pip_5160_1_126___stage___block_26_v_x[2+:2]};

_t___stage___block_2540_vnum2 = {_q___pip_5160_1_126___stage___block_26_v_z[4+:2],_q___pip_5160_1_126___stage___block_26_v_y[4+:2],_q___pip_5160_1_126___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_126___stage___block_6_inside&_w_tile[_t___stage___block_2540_vnum0+:1]&_w_tile[_t___stage___block_2540_vnum1+:1]&_w_tile[_t___stage___block_2540_vnum2+:1]) begin
// __block_2541
// __block_2543
_d___pip_5160_1_126___stage___block_6_clr = _t___stage___block_2540_tex;

_d___pip_5160_1_126___stage___block_6_dist = 222;

_d___pip_5160_1_126___stage___block_6_inside = 1;

// __block_2544
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2542
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2545
_t___block_2545_cmp_yx = _q___pip_5160_1_126___block_34_tm_y-_q___pip_5160_1_126___block_34_tm_x;

_t___block_2545_cmp_zx = _q___pip_5160_1_126___block_34_tm_z-_q___pip_5160_1_126___block_34_tm_x;

_t___block_2545_cmp_zy = _q___pip_5160_1_126___block_34_tm_z-_q___pip_5160_1_126___block_34_tm_y;

_t___block_2545_x_sel = ~_t___block_2545_cmp_yx[20+:1]&&~_t___block_2545_cmp_zx[20+:1];

_t___block_2545_y_sel = _t___block_2545_cmp_yx[20+:1]&&~_t___block_2545_cmp_zy[20+:1];

_t___block_2545_z_sel = _t___block_2545_cmp_zx[20+:1]&&_t___block_2545_cmp_zy[20+:1];

if (_t___block_2545_x_sel) begin
// __block_2546
// __block_2548
_d___pip_5160_1_126___stage___block_26_v_x = _q___pip_5160_1_126___stage___block_26_v_x+_q___pip_5160_1_126___stage___block_26_s_x;

_d___pip_5160_1_126___block_34_tm_x = _q___pip_5160_1_126___block_34_tm_x+_q___pip_5160_1_126___block_40_dt_x;

// __block_2549
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2547
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2550
if (_t___block_2545_y_sel) begin
// __block_2551
// __block_2553
_d___pip_5160_1_126___stage___block_26_v_y = _q___pip_5160_1_126___stage___block_26_v_y+_q___pip_5160_1_126___stage___block_26_s_y;

_d___pip_5160_1_126___block_34_tm_y = _q___pip_5160_1_126___block_34_tm_y+_q___pip_5160_1_126___block_40_dt_y;

// __block_2554
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2552
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2555
if (_t___block_2545_z_sel) begin
// __block_2556
// __block_2558
_d___pip_5160_1_126___stage___block_26_v_z = _q___pip_5160_1_126___stage___block_26_v_z+_q___pip_5160_1_126___stage___block_26_s_z;

_d___pip_5160_1_126___block_34_tm_z = _q___pip_5160_1_126___block_34_tm_z+_q___pip_5160_1_126___block_40_dt_z;

// __block_2559
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2557
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2560
// end of pipeline stage
_d__full_fsm___pip_5160_1_126 = 1;
_d__idx_fsm___pip_5160_1_126 = _t__stall_fsm___pip_5160_1_126 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_126 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 127
(* full_case *)
case (_q__idx_fsm___pip_5160_1_127)
1: begin
// __stage___block_2561
_t___stage___block_2561_tex = (_q___pip_5160_1_127___stage___block_26_v_x)^(_q___pip_5160_1_127___stage___block_26_v_y)^(_q___pip_5160_1_127___stage___block_26_v_z);

_t___stage___block_2561_vnum0 = {_q___pip_5160_1_127___stage___block_26_v_z[0+:2],_q___pip_5160_1_127___stage___block_26_v_y[0+:2],_q___pip_5160_1_127___stage___block_26_v_x[0+:2]};

_t___stage___block_2561_vnum1 = {_q___pip_5160_1_127___stage___block_26_v_z[2+:2],_q___pip_5160_1_127___stage___block_26_v_y[2+:2],_q___pip_5160_1_127___stage___block_26_v_x[2+:2]};

_t___stage___block_2561_vnum2 = {_q___pip_5160_1_127___stage___block_26_v_z[4+:2],_q___pip_5160_1_127___stage___block_26_v_y[4+:2],_q___pip_5160_1_127___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_127___stage___block_6_inside&_w_tile[_t___stage___block_2561_vnum0+:1]&_w_tile[_t___stage___block_2561_vnum1+:1]&_w_tile[_t___stage___block_2561_vnum2+:1]) begin
// __block_2562
// __block_2564
_d___pip_5160_1_127___stage___block_6_clr = _t___stage___block_2561_tex;

_d___pip_5160_1_127___stage___block_6_dist = 224;

_d___pip_5160_1_127___stage___block_6_inside = 1;

// __block_2565
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2563
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2566
_t___block_2566_cmp_yx = _q___pip_5160_1_127___block_34_tm_y-_q___pip_5160_1_127___block_34_tm_x;

_t___block_2566_cmp_zx = _q___pip_5160_1_127___block_34_tm_z-_q___pip_5160_1_127___block_34_tm_x;

_t___block_2566_cmp_zy = _q___pip_5160_1_127___block_34_tm_z-_q___pip_5160_1_127___block_34_tm_y;

_t___block_2566_x_sel = ~_t___block_2566_cmp_yx[20+:1]&&~_t___block_2566_cmp_zx[20+:1];

_t___block_2566_y_sel = _t___block_2566_cmp_yx[20+:1]&&~_t___block_2566_cmp_zy[20+:1];

_t___block_2566_z_sel = _t___block_2566_cmp_zx[20+:1]&&_t___block_2566_cmp_zy[20+:1];

if (_t___block_2566_x_sel) begin
// __block_2567
// __block_2569
_d___pip_5160_1_127___stage___block_26_v_x = _q___pip_5160_1_127___stage___block_26_v_x+_q___pip_5160_1_127___stage___block_26_s_x;

_d___pip_5160_1_127___block_34_tm_x = _q___pip_5160_1_127___block_34_tm_x+_q___pip_5160_1_127___block_40_dt_x;

// __block_2570
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2568
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2571
if (_t___block_2566_y_sel) begin
// __block_2572
// __block_2574
_d___pip_5160_1_127___stage___block_26_v_y = _q___pip_5160_1_127___stage___block_26_v_y+_q___pip_5160_1_127___stage___block_26_s_y;

_d___pip_5160_1_127___block_34_tm_y = _q___pip_5160_1_127___block_34_tm_y+_q___pip_5160_1_127___block_40_dt_y;

// __block_2575
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2573
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2576
if (_t___block_2566_z_sel) begin
// __block_2577
// __block_2579
_d___pip_5160_1_127___stage___block_26_v_z = _q___pip_5160_1_127___stage___block_26_v_z+_q___pip_5160_1_127___stage___block_26_s_z;

_d___pip_5160_1_127___block_34_tm_z = _q___pip_5160_1_127___block_34_tm_z+_q___pip_5160_1_127___block_40_dt_z;

// __block_2580
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2578
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2581
// end of pipeline stage
_d__full_fsm___pip_5160_1_127 = 1;
_d__idx_fsm___pip_5160_1_127 = _t__stall_fsm___pip_5160_1_127 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_127 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 128
(* full_case *)
case (_q__idx_fsm___pip_5160_1_128)
1: begin
// __stage___block_2582
_t___stage___block_2582_tex = (_q___pip_5160_1_128___stage___block_26_v_x)^(_q___pip_5160_1_128___stage___block_26_v_y)^(_q___pip_5160_1_128___stage___block_26_v_z);

_t___stage___block_2582_vnum0 = {_q___pip_5160_1_128___stage___block_26_v_z[0+:2],_q___pip_5160_1_128___stage___block_26_v_y[0+:2],_q___pip_5160_1_128___stage___block_26_v_x[0+:2]};

_t___stage___block_2582_vnum1 = {_q___pip_5160_1_128___stage___block_26_v_z[2+:2],_q___pip_5160_1_128___stage___block_26_v_y[2+:2],_q___pip_5160_1_128___stage___block_26_v_x[2+:2]};

_t___stage___block_2582_vnum2 = {_q___pip_5160_1_128___stage___block_26_v_z[4+:2],_q___pip_5160_1_128___stage___block_26_v_y[4+:2],_q___pip_5160_1_128___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_128___stage___block_6_inside&_w_tile[_t___stage___block_2582_vnum0+:1]&_w_tile[_t___stage___block_2582_vnum1+:1]&_w_tile[_t___stage___block_2582_vnum2+:1]) begin
// __block_2583
// __block_2585
_d___pip_5160_1_128___stage___block_6_clr = _t___stage___block_2582_tex;

_d___pip_5160_1_128___stage___block_6_dist = 225;

_d___pip_5160_1_128___stage___block_6_inside = 1;

// __block_2586
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2584
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2587
_t___block_2587_cmp_yx = _q___pip_5160_1_128___block_34_tm_y-_q___pip_5160_1_128___block_34_tm_x;

_t___block_2587_cmp_zx = _q___pip_5160_1_128___block_34_tm_z-_q___pip_5160_1_128___block_34_tm_x;

_t___block_2587_cmp_zy = _q___pip_5160_1_128___block_34_tm_z-_q___pip_5160_1_128___block_34_tm_y;

_t___block_2587_x_sel = ~_t___block_2587_cmp_yx[20+:1]&&~_t___block_2587_cmp_zx[20+:1];

_t___block_2587_y_sel = _t___block_2587_cmp_yx[20+:1]&&~_t___block_2587_cmp_zy[20+:1];

_t___block_2587_z_sel = _t___block_2587_cmp_zx[20+:1]&&_t___block_2587_cmp_zy[20+:1];

if (_t___block_2587_x_sel) begin
// __block_2588
// __block_2590
_d___pip_5160_1_128___stage___block_26_v_x = _q___pip_5160_1_128___stage___block_26_v_x+_q___pip_5160_1_128___stage___block_26_s_x;

_d___pip_5160_1_128___block_34_tm_x = _q___pip_5160_1_128___block_34_tm_x+_q___pip_5160_1_128___block_40_dt_x;

// __block_2591
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2589
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2592
if (_t___block_2587_y_sel) begin
// __block_2593
// __block_2595
_d___pip_5160_1_128___stage___block_26_v_y = _q___pip_5160_1_128___stage___block_26_v_y+_q___pip_5160_1_128___stage___block_26_s_y;

_d___pip_5160_1_128___block_34_tm_y = _q___pip_5160_1_128___block_34_tm_y+_q___pip_5160_1_128___block_40_dt_y;

// __block_2596
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2594
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2597
if (_t___block_2587_z_sel) begin
// __block_2598
// __block_2600
_d___pip_5160_1_128___stage___block_26_v_z = _q___pip_5160_1_128___stage___block_26_v_z+_q___pip_5160_1_128___stage___block_26_s_z;

_d___pip_5160_1_128___block_34_tm_z = _q___pip_5160_1_128___block_34_tm_z+_q___pip_5160_1_128___block_40_dt_z;

// __block_2601
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2599
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2602
// end of pipeline stage
_d__full_fsm___pip_5160_1_128 = 1;
_d__idx_fsm___pip_5160_1_128 = _t__stall_fsm___pip_5160_1_128 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_128 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 129
(* full_case *)
case (_q__idx_fsm___pip_5160_1_129)
1: begin
// __stage___block_2603
_t___stage___block_2603_tex = (_q___pip_5160_1_129___stage___block_26_v_x)^(_q___pip_5160_1_129___stage___block_26_v_y)^(_q___pip_5160_1_129___stage___block_26_v_z);

_t___stage___block_2603_vnum0 = {_q___pip_5160_1_129___stage___block_26_v_z[0+:2],_q___pip_5160_1_129___stage___block_26_v_y[0+:2],_q___pip_5160_1_129___stage___block_26_v_x[0+:2]};

_t___stage___block_2603_vnum1 = {_q___pip_5160_1_129___stage___block_26_v_z[2+:2],_q___pip_5160_1_129___stage___block_26_v_y[2+:2],_q___pip_5160_1_129___stage___block_26_v_x[2+:2]};

_t___stage___block_2603_vnum2 = {_q___pip_5160_1_129___stage___block_26_v_z[4+:2],_q___pip_5160_1_129___stage___block_26_v_y[4+:2],_q___pip_5160_1_129___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_129___stage___block_6_inside&_w_tile[_t___stage___block_2603_vnum0+:1]&_w_tile[_t___stage___block_2603_vnum1+:1]&_w_tile[_t___stage___block_2603_vnum2+:1]) begin
// __block_2604
// __block_2606
_d___pip_5160_1_129___stage___block_6_clr = _t___stage___block_2603_tex;

_d___pip_5160_1_129___stage___block_6_dist = 227;

_d___pip_5160_1_129___stage___block_6_inside = 1;

// __block_2607
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2605
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2608
_t___block_2608_cmp_yx = _q___pip_5160_1_129___block_34_tm_y-_q___pip_5160_1_129___block_34_tm_x;

_t___block_2608_cmp_zx = _q___pip_5160_1_129___block_34_tm_z-_q___pip_5160_1_129___block_34_tm_x;

_t___block_2608_cmp_zy = _q___pip_5160_1_129___block_34_tm_z-_q___pip_5160_1_129___block_34_tm_y;

_t___block_2608_x_sel = ~_t___block_2608_cmp_yx[20+:1]&&~_t___block_2608_cmp_zx[20+:1];

_t___block_2608_y_sel = _t___block_2608_cmp_yx[20+:1]&&~_t___block_2608_cmp_zy[20+:1];

_t___block_2608_z_sel = _t___block_2608_cmp_zx[20+:1]&&_t___block_2608_cmp_zy[20+:1];

if (_t___block_2608_x_sel) begin
// __block_2609
// __block_2611
_d___pip_5160_1_129___stage___block_26_v_x = _q___pip_5160_1_129___stage___block_26_v_x+_q___pip_5160_1_129___stage___block_26_s_x;

_d___pip_5160_1_129___block_34_tm_x = _q___pip_5160_1_129___block_34_tm_x+_q___pip_5160_1_129___block_40_dt_x;

// __block_2612
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2610
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2613
if (_t___block_2608_y_sel) begin
// __block_2614
// __block_2616
_d___pip_5160_1_129___stage___block_26_v_y = _q___pip_5160_1_129___stage___block_26_v_y+_q___pip_5160_1_129___stage___block_26_s_y;

_d___pip_5160_1_129___block_34_tm_y = _q___pip_5160_1_129___block_34_tm_y+_q___pip_5160_1_129___block_40_dt_y;

// __block_2617
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2615
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2618
if (_t___block_2608_z_sel) begin
// __block_2619
// __block_2621
_d___pip_5160_1_129___stage___block_26_v_z = _q___pip_5160_1_129___stage___block_26_v_z+_q___pip_5160_1_129___stage___block_26_s_z;

_d___pip_5160_1_129___block_34_tm_z = _q___pip_5160_1_129___block_34_tm_z+_q___pip_5160_1_129___block_40_dt_z;

// __block_2622
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2620
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2623
// end of pipeline stage
_d__full_fsm___pip_5160_1_129 = 1;
_d__idx_fsm___pip_5160_1_129 = _t__stall_fsm___pip_5160_1_129 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_129 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 130
(* full_case *)
case (_q__idx_fsm___pip_5160_1_130)
1: begin
// __stage___block_2624
_t___stage___block_2624_tex = (_q___pip_5160_1_130___stage___block_26_v_x)^(_q___pip_5160_1_130___stage___block_26_v_y)^(_q___pip_5160_1_130___stage___block_26_v_z);

_t___stage___block_2624_vnum0 = {_q___pip_5160_1_130___stage___block_26_v_z[0+:2],_q___pip_5160_1_130___stage___block_26_v_y[0+:2],_q___pip_5160_1_130___stage___block_26_v_x[0+:2]};

_t___stage___block_2624_vnum1 = {_q___pip_5160_1_130___stage___block_26_v_z[2+:2],_q___pip_5160_1_130___stage___block_26_v_y[2+:2],_q___pip_5160_1_130___stage___block_26_v_x[2+:2]};

_t___stage___block_2624_vnum2 = {_q___pip_5160_1_130___stage___block_26_v_z[4+:2],_q___pip_5160_1_130___stage___block_26_v_y[4+:2],_q___pip_5160_1_130___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_130___stage___block_6_inside&_w_tile[_t___stage___block_2624_vnum0+:1]&_w_tile[_t___stage___block_2624_vnum1+:1]&_w_tile[_t___stage___block_2624_vnum2+:1]) begin
// __block_2625
// __block_2627
_d___pip_5160_1_130___stage___block_6_clr = _t___stage___block_2624_tex;

_d___pip_5160_1_130___stage___block_6_dist = 229;

_d___pip_5160_1_130___stage___block_6_inside = 1;

// __block_2628
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2626
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2629
_t___block_2629_cmp_yx = _q___pip_5160_1_130___block_34_tm_y-_q___pip_5160_1_130___block_34_tm_x;

_t___block_2629_cmp_zx = _q___pip_5160_1_130___block_34_tm_z-_q___pip_5160_1_130___block_34_tm_x;

_t___block_2629_cmp_zy = _q___pip_5160_1_130___block_34_tm_z-_q___pip_5160_1_130___block_34_tm_y;

_t___block_2629_x_sel = ~_t___block_2629_cmp_yx[20+:1]&&~_t___block_2629_cmp_zx[20+:1];

_t___block_2629_y_sel = _t___block_2629_cmp_yx[20+:1]&&~_t___block_2629_cmp_zy[20+:1];

_t___block_2629_z_sel = _t___block_2629_cmp_zx[20+:1]&&_t___block_2629_cmp_zy[20+:1];

if (_t___block_2629_x_sel) begin
// __block_2630
// __block_2632
_d___pip_5160_1_130___stage___block_26_v_x = _q___pip_5160_1_130___stage___block_26_v_x+_q___pip_5160_1_130___stage___block_26_s_x;

_d___pip_5160_1_130___block_34_tm_x = _q___pip_5160_1_130___block_34_tm_x+_q___pip_5160_1_130___block_40_dt_x;

// __block_2633
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2631
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2634
if (_t___block_2629_y_sel) begin
// __block_2635
// __block_2637
_d___pip_5160_1_130___stage___block_26_v_y = _q___pip_5160_1_130___stage___block_26_v_y+_q___pip_5160_1_130___stage___block_26_s_y;

_d___pip_5160_1_130___block_34_tm_y = _q___pip_5160_1_130___block_34_tm_y+_q___pip_5160_1_130___block_40_dt_y;

// __block_2638
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2636
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2639
if (_t___block_2629_z_sel) begin
// __block_2640
// __block_2642
_d___pip_5160_1_130___stage___block_26_v_z = _q___pip_5160_1_130___stage___block_26_v_z+_q___pip_5160_1_130___stage___block_26_s_z;

_d___pip_5160_1_130___block_34_tm_z = _q___pip_5160_1_130___block_34_tm_z+_q___pip_5160_1_130___block_40_dt_z;

// __block_2643
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2641
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2644
// end of pipeline stage
_d__full_fsm___pip_5160_1_130 = 1;
_d__idx_fsm___pip_5160_1_130 = _t__stall_fsm___pip_5160_1_130 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_130 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 131
(* full_case *)
case (_q__idx_fsm___pip_5160_1_131)
1: begin
// __stage___block_2645
_t___stage___block_2645_tex = (_q___pip_5160_1_131___stage___block_26_v_x)^(_q___pip_5160_1_131___stage___block_26_v_y)^(_q___pip_5160_1_131___stage___block_26_v_z);

_t___stage___block_2645_vnum0 = {_q___pip_5160_1_131___stage___block_26_v_z[0+:2],_q___pip_5160_1_131___stage___block_26_v_y[0+:2],_q___pip_5160_1_131___stage___block_26_v_x[0+:2]};

_t___stage___block_2645_vnum1 = {_q___pip_5160_1_131___stage___block_26_v_z[2+:2],_q___pip_5160_1_131___stage___block_26_v_y[2+:2],_q___pip_5160_1_131___stage___block_26_v_x[2+:2]};

_t___stage___block_2645_vnum2 = {_q___pip_5160_1_131___stage___block_26_v_z[4+:2],_q___pip_5160_1_131___stage___block_26_v_y[4+:2],_q___pip_5160_1_131___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_131___stage___block_6_inside&_w_tile[_t___stage___block_2645_vnum0+:1]&_w_tile[_t___stage___block_2645_vnum1+:1]&_w_tile[_t___stage___block_2645_vnum2+:1]) begin
// __block_2646
// __block_2648
_d___pip_5160_1_131___stage___block_6_clr = _t___stage___block_2645_tex;

_d___pip_5160_1_131___stage___block_6_dist = 231;

_d___pip_5160_1_131___stage___block_6_inside = 1;

// __block_2649
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2647
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2650
_t___block_2650_cmp_yx = _q___pip_5160_1_131___block_34_tm_y-_q___pip_5160_1_131___block_34_tm_x;

_t___block_2650_cmp_zx = _q___pip_5160_1_131___block_34_tm_z-_q___pip_5160_1_131___block_34_tm_x;

_t___block_2650_cmp_zy = _q___pip_5160_1_131___block_34_tm_z-_q___pip_5160_1_131___block_34_tm_y;

_t___block_2650_x_sel = ~_t___block_2650_cmp_yx[20+:1]&&~_t___block_2650_cmp_zx[20+:1];

_t___block_2650_y_sel = _t___block_2650_cmp_yx[20+:1]&&~_t___block_2650_cmp_zy[20+:1];

_t___block_2650_z_sel = _t___block_2650_cmp_zx[20+:1]&&_t___block_2650_cmp_zy[20+:1];

if (_t___block_2650_x_sel) begin
// __block_2651
// __block_2653
_d___pip_5160_1_131___stage___block_26_v_x = _q___pip_5160_1_131___stage___block_26_v_x+_q___pip_5160_1_131___stage___block_26_s_x;

_d___pip_5160_1_131___block_34_tm_x = _q___pip_5160_1_131___block_34_tm_x+_q___pip_5160_1_131___block_40_dt_x;

// __block_2654
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2652
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2655
if (_t___block_2650_y_sel) begin
// __block_2656
// __block_2658
_d___pip_5160_1_131___stage___block_26_v_y = _q___pip_5160_1_131___stage___block_26_v_y+_q___pip_5160_1_131___stage___block_26_s_y;

_d___pip_5160_1_131___block_34_tm_y = _q___pip_5160_1_131___block_34_tm_y+_q___pip_5160_1_131___block_40_dt_y;

// __block_2659
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2657
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2660
if (_t___block_2650_z_sel) begin
// __block_2661
// __block_2663
_d___pip_5160_1_131___stage___block_26_v_z = _q___pip_5160_1_131___stage___block_26_v_z+_q___pip_5160_1_131___stage___block_26_s_z;

_d___pip_5160_1_131___block_34_tm_z = _q___pip_5160_1_131___block_34_tm_z+_q___pip_5160_1_131___block_40_dt_z;

// __block_2664
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2662
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2665
// end of pipeline stage
_d__full_fsm___pip_5160_1_131 = 1;
_d__idx_fsm___pip_5160_1_131 = _t__stall_fsm___pip_5160_1_131 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_131 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 132
(* full_case *)
case (_q__idx_fsm___pip_5160_1_132)
1: begin
// __stage___block_2666
_t___stage___block_2666_tex = (_q___pip_5160_1_132___stage___block_26_v_x)^(_q___pip_5160_1_132___stage___block_26_v_y)^(_q___pip_5160_1_132___stage___block_26_v_z);

_t___stage___block_2666_vnum0 = {_q___pip_5160_1_132___stage___block_26_v_z[0+:2],_q___pip_5160_1_132___stage___block_26_v_y[0+:2],_q___pip_5160_1_132___stage___block_26_v_x[0+:2]};

_t___stage___block_2666_vnum1 = {_q___pip_5160_1_132___stage___block_26_v_z[2+:2],_q___pip_5160_1_132___stage___block_26_v_y[2+:2],_q___pip_5160_1_132___stage___block_26_v_x[2+:2]};

_t___stage___block_2666_vnum2 = {_q___pip_5160_1_132___stage___block_26_v_z[4+:2],_q___pip_5160_1_132___stage___block_26_v_y[4+:2],_q___pip_5160_1_132___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_132___stage___block_6_inside&_w_tile[_t___stage___block_2666_vnum0+:1]&_w_tile[_t___stage___block_2666_vnum1+:1]&_w_tile[_t___stage___block_2666_vnum2+:1]) begin
// __block_2667
// __block_2669
_d___pip_5160_1_132___stage___block_6_clr = _t___stage___block_2666_tex;

_d___pip_5160_1_132___stage___block_6_dist = 233;

_d___pip_5160_1_132___stage___block_6_inside = 1;

// __block_2670
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2668
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2671
_t___block_2671_cmp_yx = _q___pip_5160_1_132___block_34_tm_y-_q___pip_5160_1_132___block_34_tm_x;

_t___block_2671_cmp_zx = _q___pip_5160_1_132___block_34_tm_z-_q___pip_5160_1_132___block_34_tm_x;

_t___block_2671_cmp_zy = _q___pip_5160_1_132___block_34_tm_z-_q___pip_5160_1_132___block_34_tm_y;

_t___block_2671_x_sel = ~_t___block_2671_cmp_yx[20+:1]&&~_t___block_2671_cmp_zx[20+:1];

_t___block_2671_y_sel = _t___block_2671_cmp_yx[20+:1]&&~_t___block_2671_cmp_zy[20+:1];

_t___block_2671_z_sel = _t___block_2671_cmp_zx[20+:1]&&_t___block_2671_cmp_zy[20+:1];

if (_t___block_2671_x_sel) begin
// __block_2672
// __block_2674
_d___pip_5160_1_132___stage___block_26_v_x = _q___pip_5160_1_132___stage___block_26_v_x+_q___pip_5160_1_132___stage___block_26_s_x;

_d___pip_5160_1_132___block_34_tm_x = _q___pip_5160_1_132___block_34_tm_x+_q___pip_5160_1_132___block_40_dt_x;

// __block_2675
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2673
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2676
if (_t___block_2671_y_sel) begin
// __block_2677
// __block_2679
_d___pip_5160_1_132___stage___block_26_v_y = _q___pip_5160_1_132___stage___block_26_v_y+_q___pip_5160_1_132___stage___block_26_s_y;

_d___pip_5160_1_132___block_34_tm_y = _q___pip_5160_1_132___block_34_tm_y+_q___pip_5160_1_132___block_40_dt_y;

// __block_2680
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2678
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2681
if (_t___block_2671_z_sel) begin
// __block_2682
// __block_2684
_d___pip_5160_1_132___stage___block_26_v_z = _q___pip_5160_1_132___stage___block_26_v_z+_q___pip_5160_1_132___stage___block_26_s_z;

_d___pip_5160_1_132___block_34_tm_z = _q___pip_5160_1_132___block_34_tm_z+_q___pip_5160_1_132___block_40_dt_z;

// __block_2685
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2683
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2686
// end of pipeline stage
_d__full_fsm___pip_5160_1_132 = 1;
_d__idx_fsm___pip_5160_1_132 = _t__stall_fsm___pip_5160_1_132 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_132 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 133
(* full_case *)
case (_q__idx_fsm___pip_5160_1_133)
1: begin
// __stage___block_2687
_t___stage___block_2687_tex = (_q___pip_5160_1_133___stage___block_26_v_x)^(_q___pip_5160_1_133___stage___block_26_v_y)^(_q___pip_5160_1_133___stage___block_26_v_z);

_t___stage___block_2687_vnum0 = {_q___pip_5160_1_133___stage___block_26_v_z[0+:2],_q___pip_5160_1_133___stage___block_26_v_y[0+:2],_q___pip_5160_1_133___stage___block_26_v_x[0+:2]};

_t___stage___block_2687_vnum1 = {_q___pip_5160_1_133___stage___block_26_v_z[2+:2],_q___pip_5160_1_133___stage___block_26_v_y[2+:2],_q___pip_5160_1_133___stage___block_26_v_x[2+:2]};

_t___stage___block_2687_vnum2 = {_q___pip_5160_1_133___stage___block_26_v_z[4+:2],_q___pip_5160_1_133___stage___block_26_v_y[4+:2],_q___pip_5160_1_133___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_133___stage___block_6_inside&_w_tile[_t___stage___block_2687_vnum0+:1]&_w_tile[_t___stage___block_2687_vnum1+:1]&_w_tile[_t___stage___block_2687_vnum2+:1]) begin
// __block_2688
// __block_2690
_d___pip_5160_1_133___stage___block_6_clr = _t___stage___block_2687_tex;

_d___pip_5160_1_133___stage___block_6_dist = 235;

_d___pip_5160_1_133___stage___block_6_inside = 1;

// __block_2691
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2689
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2692
_t___block_2692_cmp_yx = _q___pip_5160_1_133___block_34_tm_y-_q___pip_5160_1_133___block_34_tm_x;

_t___block_2692_cmp_zx = _q___pip_5160_1_133___block_34_tm_z-_q___pip_5160_1_133___block_34_tm_x;

_t___block_2692_cmp_zy = _q___pip_5160_1_133___block_34_tm_z-_q___pip_5160_1_133___block_34_tm_y;

_t___block_2692_x_sel = ~_t___block_2692_cmp_yx[20+:1]&&~_t___block_2692_cmp_zx[20+:1];

_t___block_2692_y_sel = _t___block_2692_cmp_yx[20+:1]&&~_t___block_2692_cmp_zy[20+:1];

_t___block_2692_z_sel = _t___block_2692_cmp_zx[20+:1]&&_t___block_2692_cmp_zy[20+:1];

if (_t___block_2692_x_sel) begin
// __block_2693
// __block_2695
_d___pip_5160_1_133___stage___block_26_v_x = _q___pip_5160_1_133___stage___block_26_v_x+_q___pip_5160_1_133___stage___block_26_s_x;

_d___pip_5160_1_133___block_34_tm_x = _q___pip_5160_1_133___block_34_tm_x+_q___pip_5160_1_133___block_40_dt_x;

// __block_2696
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2694
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2697
if (_t___block_2692_y_sel) begin
// __block_2698
// __block_2700
_d___pip_5160_1_133___stage___block_26_v_y = _q___pip_5160_1_133___stage___block_26_v_y+_q___pip_5160_1_133___stage___block_26_s_y;

_d___pip_5160_1_133___block_34_tm_y = _q___pip_5160_1_133___block_34_tm_y+_q___pip_5160_1_133___block_40_dt_y;

// __block_2701
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2699
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2702
if (_t___block_2692_z_sel) begin
// __block_2703
// __block_2705
_d___pip_5160_1_133___stage___block_26_v_z = _q___pip_5160_1_133___stage___block_26_v_z+_q___pip_5160_1_133___stage___block_26_s_z;

_d___pip_5160_1_133___block_34_tm_z = _q___pip_5160_1_133___block_34_tm_z+_q___pip_5160_1_133___block_40_dt_z;

// __block_2706
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2704
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2707
// end of pipeline stage
_d__full_fsm___pip_5160_1_133 = 1;
_d__idx_fsm___pip_5160_1_133 = _t__stall_fsm___pip_5160_1_133 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_133 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 134
(* full_case *)
case (_q__idx_fsm___pip_5160_1_134)
1: begin
// __stage___block_2708
_t___stage___block_2708_tex = (_q___pip_5160_1_134___stage___block_26_v_x)^(_q___pip_5160_1_134___stage___block_26_v_y)^(_q___pip_5160_1_134___stage___block_26_v_z);

_t___stage___block_2708_vnum0 = {_q___pip_5160_1_134___stage___block_26_v_z[0+:2],_q___pip_5160_1_134___stage___block_26_v_y[0+:2],_q___pip_5160_1_134___stage___block_26_v_x[0+:2]};

_t___stage___block_2708_vnum1 = {_q___pip_5160_1_134___stage___block_26_v_z[2+:2],_q___pip_5160_1_134___stage___block_26_v_y[2+:2],_q___pip_5160_1_134___stage___block_26_v_x[2+:2]};

_t___stage___block_2708_vnum2 = {_q___pip_5160_1_134___stage___block_26_v_z[4+:2],_q___pip_5160_1_134___stage___block_26_v_y[4+:2],_q___pip_5160_1_134___stage___block_26_v_x[4+:2]};

if (~_q___pip_5160_1_134___stage___block_6_inside&_w_tile[_t___stage___block_2708_vnum0+:1]&_w_tile[_t___stage___block_2708_vnum1+:1]&_w_tile[_t___stage___block_2708_vnum2+:1]) begin
// __block_2709
// __block_2711
_d___pip_5160_1_134___stage___block_6_clr = _t___stage___block_2708_tex;

_d___pip_5160_1_134___stage___block_6_dist = 237;

_d___pip_5160_1_134___stage___block_6_inside = 1;

// __block_2712
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2710
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2713
_t___block_2713_cmp_yx = _q___pip_5160_1_134___block_34_tm_y-_q___pip_5160_1_134___block_34_tm_x;

_t___block_2713_cmp_zx = _q___pip_5160_1_134___block_34_tm_z-_q___pip_5160_1_134___block_34_tm_x;

_t___block_2713_cmp_zy = _q___pip_5160_1_134___block_34_tm_z-_q___pip_5160_1_134___block_34_tm_y;

_t___block_2713_x_sel = ~_t___block_2713_cmp_yx[20+:1]&&~_t___block_2713_cmp_zx[20+:1];

_t___block_2713_y_sel = _t___block_2713_cmp_yx[20+:1]&&~_t___block_2713_cmp_zy[20+:1];

_t___block_2713_z_sel = _t___block_2713_cmp_zx[20+:1]&&_t___block_2713_cmp_zy[20+:1];

if (_t___block_2713_x_sel) begin
// __block_2714
// __block_2716
_d___pip_5160_1_134___stage___block_26_v_x = _q___pip_5160_1_134___stage___block_26_v_x+_q___pip_5160_1_134___stage___block_26_s_x;

_d___pip_5160_1_134___block_34_tm_x = _q___pip_5160_1_134___block_34_tm_x+_q___pip_5160_1_134___block_40_dt_x;

// __block_2717
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2715
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2718
if (_t___block_2713_y_sel) begin
// __block_2719
// __block_2721
_d___pip_5160_1_134___stage___block_26_v_y = _q___pip_5160_1_134___stage___block_26_v_y+_q___pip_5160_1_134___stage___block_26_s_y;

_d___pip_5160_1_134___block_34_tm_y = _q___pip_5160_1_134___block_34_tm_y+_q___pip_5160_1_134___block_40_dt_y;

// __block_2722
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2720
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2723
if (_t___block_2713_z_sel) begin
// __block_2724
// __block_2726
_d___pip_5160_1_134___stage___block_26_v_z = _q___pip_5160_1_134___stage___block_26_v_z+_q___pip_5160_1_134___stage___block_26_s_z;

_d___pip_5160_1_134___block_34_tm_z = _q___pip_5160_1_134___block_34_tm_z+_q___pip_5160_1_134___block_40_dt_z;

// __block_2727
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end else begin
// __block_2725
_t__1stdisable_fsm___pip_5160_1_0 = 1;
end
// 'after'
// __block_2728
// end of pipeline stage
_d__full_fsm___pip_5160_1_134 = 1;
_d__idx_fsm___pip_5160_1_134 = _t__stall_fsm___pip_5160_1_134 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_134 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// -------- stage 135
(* full_case *)
case (_q__idx_fsm___pip_5160_1_135)
1: begin
// __stage___block_2729
_t___stage___block_2729_fog = _q___pip_5160_1_135___stage___block_6_dist;

_t___stage___block_2729_light = 239-_t___stage___block_2729_fog;

// __block_2730_mul_8_8
_t___stage___block_2729_shade = _t___stage___block_2729_light*_q___pip_5160_1_135___stage___block_6_clr;

// __block_2731
_t___block_2731_clr_r = (_t___stage___block_2729_shade[7+:8])+_t___stage___block_2729_fog;

_t___block_2731_clr_g = (_t___stage___block_2729_shade[7+:8])+_t___stage___block_2729_fog;

_t___block_2731_clr_b = (_t___stage___block_2729_shade[8+:8])+_t___stage___block_2729_fog;

// end of pipeline stage
_d__full_fsm___pip_5160_1_135 = 1;
_d__idx_fsm___pip_5160_1_135 = _t__stall_fsm___pip_5160_1_135 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_135 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
if (_q__idx_fsm___pip_5160_1_135 == 1  ) begin
_d___pip_5160_1_135___block_2731_clr_r = _t___block_2731_clr_r;
end else begin
_d___pip_5160_1_135___block_2731_clr_r = _q___pip_5160_1_135___block_2731_clr_r;
end
if (_q__idx_fsm___pip_5160_1_135 == 1  ) begin
_d___pip_5160_1_135___block_2731_clr_g = _t___block_2731_clr_g;
end else begin
_d___pip_5160_1_135___block_2731_clr_g = _q___pip_5160_1_135___block_2731_clr_g;
end
if (_q__idx_fsm___pip_5160_1_135 == 1  ) begin
_d___pip_5160_1_135___block_2731_clr_b = _t___block_2731_clr_b;
end else begin
_d___pip_5160_1_135___block_2731_clr_b = _q___pip_5160_1_135___block_2731_clr_b;
end
// -------- stage 136
(* full_case *)
case (_q__idx_fsm___pip_5160_1_136)
1: begin
// __stage___block_2732
_d_pix_r = _q___pip_5160_1_136___block_2731_clr_r;

_d_pix_g = _q___pip_5160_1_136___block_2731_clr_g;

_d_pix_b = _q___pip_5160_1_136___block_2731_clr_b;

if (in_pix_x==0&&in_pix_y==0) begin
// __block_2733
// __block_2735
_d_frame = (_q_frame-1);

// __block_2736
end else begin
// __block_2734
end
// 'after'
// __block_2737
// end of last pipeline stage
_d__full_fsm___pip_5160_1_136 = 1;
_d__idx_fsm___pip_5160_1_136 = _t__stall_fsm___pip_5160_1_136 ? 1 : 0;
end
0: begin 
end
default: begin 
_d__idx_fsm___pip_5160_1_136 = {1{1'bx}};
`ifdef FORMAL
assume(0);
`endif
 end
endcase
// --- trickling
// ===================
// _always_post
// pipeline stage triggers
if ( (_ready_fsm___pip_5160_1_136)   && (_d__full_fsm___pip_5160_1_135)   && (!_t__stall_fsm___pip_5160_1_135)   && (!_t__stall_fsm___pip_5160_1_136)   ) begin
   _d__idx_fsm___pip_5160_1_136 = 1;
   _d__full_fsm___pip_5160_1_135 = 0;
end
if ( (_ready_fsm___pip_5160_1_135)   && (_d__full_fsm___pip_5160_1_134)   && (!_t__stall_fsm___pip_5160_1_134)   && (!_d__full_fsm___pip_5160_1_135)   && (!_t__stall_fsm___pip_5160_1_135)   ) begin
   _d__idx_fsm___pip_5160_1_135 = 1;
   _d__full_fsm___pip_5160_1_134 = 0;
end
if ( (_ready_fsm___pip_5160_1_134)   && (_d__full_fsm___pip_5160_1_133)   && (!_t__stall_fsm___pip_5160_1_133)   && (!_d__full_fsm___pip_5160_1_134)   && (!_t__stall_fsm___pip_5160_1_134)   ) begin
   _d__idx_fsm___pip_5160_1_134 = 1;
   _d__full_fsm___pip_5160_1_133 = 0;
end
if ( (_ready_fsm___pip_5160_1_133)   && (_d__full_fsm___pip_5160_1_132)   && (!_t__stall_fsm___pip_5160_1_132)   && (!_d__full_fsm___pip_5160_1_133)   && (!_t__stall_fsm___pip_5160_1_133)   ) begin
   _d__idx_fsm___pip_5160_1_133 = 1;
   _d__full_fsm___pip_5160_1_132 = 0;
end
if ( (_ready_fsm___pip_5160_1_132)   && (_d__full_fsm___pip_5160_1_131)   && (!_t__stall_fsm___pip_5160_1_131)   && (!_d__full_fsm___pip_5160_1_132)   && (!_t__stall_fsm___pip_5160_1_132)   ) begin
   _d__idx_fsm___pip_5160_1_132 = 1;
   _d__full_fsm___pip_5160_1_131 = 0;
end
if ( (_ready_fsm___pip_5160_1_131)   && (_d__full_fsm___pip_5160_1_130)   && (!_t__stall_fsm___pip_5160_1_130)   && (!_d__full_fsm___pip_5160_1_131)   && (!_t__stall_fsm___pip_5160_1_131)   ) begin
   _d__idx_fsm___pip_5160_1_131 = 1;
   _d__full_fsm___pip_5160_1_130 = 0;
end
if ( (_ready_fsm___pip_5160_1_130)   && (_d__full_fsm___pip_5160_1_129)   && (!_t__stall_fsm___pip_5160_1_129)   && (!_d__full_fsm___pip_5160_1_130)   && (!_t__stall_fsm___pip_5160_1_130)   ) begin
   _d__idx_fsm___pip_5160_1_130 = 1;
   _d__full_fsm___pip_5160_1_129 = 0;
end
if ( (_ready_fsm___pip_5160_1_129)   && (_d__full_fsm___pip_5160_1_128)   && (!_t__stall_fsm___pip_5160_1_128)   && (!_d__full_fsm___pip_5160_1_129)   && (!_t__stall_fsm___pip_5160_1_129)   ) begin
   _d__idx_fsm___pip_5160_1_129 = 1;
   _d__full_fsm___pip_5160_1_128 = 0;
end
if ( (_ready_fsm___pip_5160_1_128)   && (_d__full_fsm___pip_5160_1_127)   && (!_t__stall_fsm___pip_5160_1_127)   && (!_d__full_fsm___pip_5160_1_128)   && (!_t__stall_fsm___pip_5160_1_128)   ) begin
   _d__idx_fsm___pip_5160_1_128 = 1;
   _d__full_fsm___pip_5160_1_127 = 0;
end
if ( (_ready_fsm___pip_5160_1_127)   && (_d__full_fsm___pip_5160_1_126)   && (!_t__stall_fsm___pip_5160_1_126)   && (!_d__full_fsm___pip_5160_1_127)   && (!_t__stall_fsm___pip_5160_1_127)   ) begin
   _d__idx_fsm___pip_5160_1_127 = 1;
   _d__full_fsm___pip_5160_1_126 = 0;
end
if ( (_ready_fsm___pip_5160_1_126)   && (_d__full_fsm___pip_5160_1_125)   && (!_t__stall_fsm___pip_5160_1_125)   && (!_d__full_fsm___pip_5160_1_126)   && (!_t__stall_fsm___pip_5160_1_126)   ) begin
   _d__idx_fsm___pip_5160_1_126 = 1;
   _d__full_fsm___pip_5160_1_125 = 0;
end
if ( (_ready_fsm___pip_5160_1_125)   && (_d__full_fsm___pip_5160_1_124)   && (!_t__stall_fsm___pip_5160_1_124)   && (!_d__full_fsm___pip_5160_1_125)   && (!_t__stall_fsm___pip_5160_1_125)   ) begin
   _d__idx_fsm___pip_5160_1_125 = 1;
   _d__full_fsm___pip_5160_1_124 = 0;
end
if ( (_ready_fsm___pip_5160_1_124)   && (_d__full_fsm___pip_5160_1_123)   && (!_t__stall_fsm___pip_5160_1_123)   && (!_d__full_fsm___pip_5160_1_124)   && (!_t__stall_fsm___pip_5160_1_124)   ) begin
   _d__idx_fsm___pip_5160_1_124 = 1;
   _d__full_fsm___pip_5160_1_123 = 0;
end
if ( (_ready_fsm___pip_5160_1_123)   && (_d__full_fsm___pip_5160_1_122)   && (!_t__stall_fsm___pip_5160_1_122)   && (!_d__full_fsm___pip_5160_1_123)   && (!_t__stall_fsm___pip_5160_1_123)   ) begin
   _d__idx_fsm___pip_5160_1_123 = 1;
   _d__full_fsm___pip_5160_1_122 = 0;
end
if ( (_ready_fsm___pip_5160_1_122)   && (_d__full_fsm___pip_5160_1_121)   && (!_t__stall_fsm___pip_5160_1_121)   && (!_d__full_fsm___pip_5160_1_122)   && (!_t__stall_fsm___pip_5160_1_122)   ) begin
   _d__idx_fsm___pip_5160_1_122 = 1;
   _d__full_fsm___pip_5160_1_121 = 0;
end
if ( (_ready_fsm___pip_5160_1_121)   && (_d__full_fsm___pip_5160_1_120)   && (!_t__stall_fsm___pip_5160_1_120)   && (!_d__full_fsm___pip_5160_1_121)   && (!_t__stall_fsm___pip_5160_1_121)   ) begin
   _d__idx_fsm___pip_5160_1_121 = 1;
   _d__full_fsm___pip_5160_1_120 = 0;
end
if ( (_ready_fsm___pip_5160_1_120)   && (_d__full_fsm___pip_5160_1_119)   && (!_t__stall_fsm___pip_5160_1_119)   && (!_d__full_fsm___pip_5160_1_120)   && (!_t__stall_fsm___pip_5160_1_120)   ) begin
   _d__idx_fsm___pip_5160_1_120 = 1;
   _d__full_fsm___pip_5160_1_119 = 0;
end
if ( (_ready_fsm___pip_5160_1_119)   && (_d__full_fsm___pip_5160_1_118)   && (!_t__stall_fsm___pip_5160_1_118)   && (!_d__full_fsm___pip_5160_1_119)   && (!_t__stall_fsm___pip_5160_1_119)   ) begin
   _d__idx_fsm___pip_5160_1_119 = 1;
   _d__full_fsm___pip_5160_1_118 = 0;
end
if ( (_ready_fsm___pip_5160_1_118)   && (_d__full_fsm___pip_5160_1_117)   && (!_t__stall_fsm___pip_5160_1_117)   && (!_d__full_fsm___pip_5160_1_118)   && (!_t__stall_fsm___pip_5160_1_118)   ) begin
   _d__idx_fsm___pip_5160_1_118 = 1;
   _d__full_fsm___pip_5160_1_117 = 0;
end
if ( (_ready_fsm___pip_5160_1_117)   && (_d__full_fsm___pip_5160_1_116)   && (!_t__stall_fsm___pip_5160_1_116)   && (!_d__full_fsm___pip_5160_1_117)   && (!_t__stall_fsm___pip_5160_1_117)   ) begin
   _d__idx_fsm___pip_5160_1_117 = 1;
   _d__full_fsm___pip_5160_1_116 = 0;
end
if ( (_ready_fsm___pip_5160_1_116)   && (_d__full_fsm___pip_5160_1_115)   && (!_t__stall_fsm___pip_5160_1_115)   && (!_d__full_fsm___pip_5160_1_116)   && (!_t__stall_fsm___pip_5160_1_116)   ) begin
   _d__idx_fsm___pip_5160_1_116 = 1;
   _d__full_fsm___pip_5160_1_115 = 0;
end
if ( (_ready_fsm___pip_5160_1_115)   && (_d__full_fsm___pip_5160_1_114)   && (!_t__stall_fsm___pip_5160_1_114)   && (!_d__full_fsm___pip_5160_1_115)   && (!_t__stall_fsm___pip_5160_1_115)   ) begin
   _d__idx_fsm___pip_5160_1_115 = 1;
   _d__full_fsm___pip_5160_1_114 = 0;
end
if ( (_ready_fsm___pip_5160_1_114)   && (_d__full_fsm___pip_5160_1_113)   && (!_t__stall_fsm___pip_5160_1_113)   && (!_d__full_fsm___pip_5160_1_114)   && (!_t__stall_fsm___pip_5160_1_114)   ) begin
   _d__idx_fsm___pip_5160_1_114 = 1;
   _d__full_fsm___pip_5160_1_113 = 0;
end
if ( (_ready_fsm___pip_5160_1_113)   && (_d__full_fsm___pip_5160_1_112)   && (!_t__stall_fsm___pip_5160_1_112)   && (!_d__full_fsm___pip_5160_1_113)   && (!_t__stall_fsm___pip_5160_1_113)   ) begin
   _d__idx_fsm___pip_5160_1_113 = 1;
   _d__full_fsm___pip_5160_1_112 = 0;
end
if ( (_ready_fsm___pip_5160_1_112)   && (_d__full_fsm___pip_5160_1_111)   && (!_t__stall_fsm___pip_5160_1_111)   && (!_d__full_fsm___pip_5160_1_112)   && (!_t__stall_fsm___pip_5160_1_112)   ) begin
   _d__idx_fsm___pip_5160_1_112 = 1;
   _d__full_fsm___pip_5160_1_111 = 0;
end
if ( (_ready_fsm___pip_5160_1_111)   && (_d__full_fsm___pip_5160_1_110)   && (!_t__stall_fsm___pip_5160_1_110)   && (!_d__full_fsm___pip_5160_1_111)   && (!_t__stall_fsm___pip_5160_1_111)   ) begin
   _d__idx_fsm___pip_5160_1_111 = 1;
   _d__full_fsm___pip_5160_1_110 = 0;
end
if ( (_ready_fsm___pip_5160_1_110)   && (_d__full_fsm___pip_5160_1_109)   && (!_t__stall_fsm___pip_5160_1_109)   && (!_d__full_fsm___pip_5160_1_110)   && (!_t__stall_fsm___pip_5160_1_110)   ) begin
   _d__idx_fsm___pip_5160_1_110 = 1;
   _d__full_fsm___pip_5160_1_109 = 0;
end
if ( (_ready_fsm___pip_5160_1_109)   && (_d__full_fsm___pip_5160_1_108)   && (!_t__stall_fsm___pip_5160_1_108)   && (!_d__full_fsm___pip_5160_1_109)   && (!_t__stall_fsm___pip_5160_1_109)   ) begin
   _d__idx_fsm___pip_5160_1_109 = 1;
   _d__full_fsm___pip_5160_1_108 = 0;
end
if ( (_ready_fsm___pip_5160_1_108)   && (_d__full_fsm___pip_5160_1_107)   && (!_t__stall_fsm___pip_5160_1_107)   && (!_d__full_fsm___pip_5160_1_108)   && (!_t__stall_fsm___pip_5160_1_108)   ) begin
   _d__idx_fsm___pip_5160_1_108 = 1;
   _d__full_fsm___pip_5160_1_107 = 0;
end
if ( (_ready_fsm___pip_5160_1_107)   && (_d__full_fsm___pip_5160_1_106)   && (!_t__stall_fsm___pip_5160_1_106)   && (!_d__full_fsm___pip_5160_1_107)   && (!_t__stall_fsm___pip_5160_1_107)   ) begin
   _d__idx_fsm___pip_5160_1_107 = 1;
   _d__full_fsm___pip_5160_1_106 = 0;
end
if ( (_ready_fsm___pip_5160_1_106)   && (_d__full_fsm___pip_5160_1_105)   && (!_t__stall_fsm___pip_5160_1_105)   && (!_d__full_fsm___pip_5160_1_106)   && (!_t__stall_fsm___pip_5160_1_106)   ) begin
   _d__idx_fsm___pip_5160_1_106 = 1;
   _d__full_fsm___pip_5160_1_105 = 0;
end
if ( (_ready_fsm___pip_5160_1_105)   && (_d__full_fsm___pip_5160_1_104)   && (!_t__stall_fsm___pip_5160_1_104)   && (!_d__full_fsm___pip_5160_1_105)   && (!_t__stall_fsm___pip_5160_1_105)   ) begin
   _d__idx_fsm___pip_5160_1_105 = 1;
   _d__full_fsm___pip_5160_1_104 = 0;
end
if ( (_ready_fsm___pip_5160_1_104)   && (_d__full_fsm___pip_5160_1_103)   && (!_t__stall_fsm___pip_5160_1_103)   && (!_d__full_fsm___pip_5160_1_104)   && (!_t__stall_fsm___pip_5160_1_104)   ) begin
   _d__idx_fsm___pip_5160_1_104 = 1;
   _d__full_fsm___pip_5160_1_103 = 0;
end
if ( (_ready_fsm___pip_5160_1_103)   && (_d__full_fsm___pip_5160_1_102)   && (!_t__stall_fsm___pip_5160_1_102)   && (!_d__full_fsm___pip_5160_1_103)   && (!_t__stall_fsm___pip_5160_1_103)   ) begin
   _d__idx_fsm___pip_5160_1_103 = 1;
   _d__full_fsm___pip_5160_1_102 = 0;
end
if ( (_ready_fsm___pip_5160_1_102)   && (_d__full_fsm___pip_5160_1_101)   && (!_t__stall_fsm___pip_5160_1_101)   && (!_d__full_fsm___pip_5160_1_102)   && (!_t__stall_fsm___pip_5160_1_102)   ) begin
   _d__idx_fsm___pip_5160_1_102 = 1;
   _d__full_fsm___pip_5160_1_101 = 0;
end
if ( (_ready_fsm___pip_5160_1_101)   && (_d__full_fsm___pip_5160_1_100)   && (!_t__stall_fsm___pip_5160_1_100)   && (!_d__full_fsm___pip_5160_1_101)   && (!_t__stall_fsm___pip_5160_1_101)   ) begin
   _d__idx_fsm___pip_5160_1_101 = 1;
   _d__full_fsm___pip_5160_1_100 = 0;
end
if ( (_ready_fsm___pip_5160_1_100)   && (_d__full_fsm___pip_5160_1_99)   && (!_t__stall_fsm___pip_5160_1_99)   && (!_d__full_fsm___pip_5160_1_100)   && (!_t__stall_fsm___pip_5160_1_100)   ) begin
   _d__idx_fsm___pip_5160_1_100 = 1;
   _d__full_fsm___pip_5160_1_99 = 0;
end
if ( (_ready_fsm___pip_5160_1_99)   && (_d__full_fsm___pip_5160_1_98)   && (!_t__stall_fsm___pip_5160_1_98)   && (!_d__full_fsm___pip_5160_1_99)   && (!_t__stall_fsm___pip_5160_1_99)   ) begin
   _d__idx_fsm___pip_5160_1_99 = 1;
   _d__full_fsm___pip_5160_1_98 = 0;
end
if ( (_ready_fsm___pip_5160_1_98)   && (_d__full_fsm___pip_5160_1_97)   && (!_t__stall_fsm___pip_5160_1_97)   && (!_d__full_fsm___pip_5160_1_98)   && (!_t__stall_fsm___pip_5160_1_98)   ) begin
   _d__idx_fsm___pip_5160_1_98 = 1;
   _d__full_fsm___pip_5160_1_97 = 0;
end
if ( (_ready_fsm___pip_5160_1_97)   && (_d__full_fsm___pip_5160_1_96)   && (!_t__stall_fsm___pip_5160_1_96)   && (!_d__full_fsm___pip_5160_1_97)   && (!_t__stall_fsm___pip_5160_1_97)   ) begin
   _d__idx_fsm___pip_5160_1_97 = 1;
   _d__full_fsm___pip_5160_1_96 = 0;
end
if ( (_ready_fsm___pip_5160_1_96)   && (_d__full_fsm___pip_5160_1_95)   && (!_t__stall_fsm___pip_5160_1_95)   && (!_d__full_fsm___pip_5160_1_96)   && (!_t__stall_fsm___pip_5160_1_96)   ) begin
   _d__idx_fsm___pip_5160_1_96 = 1;
   _d__full_fsm___pip_5160_1_95 = 0;
end
if ( (_ready_fsm___pip_5160_1_95)   && (_d__full_fsm___pip_5160_1_94)   && (!_t__stall_fsm___pip_5160_1_94)   && (!_d__full_fsm___pip_5160_1_95)   && (!_t__stall_fsm___pip_5160_1_95)   ) begin
   _d__idx_fsm___pip_5160_1_95 = 1;
   _d__full_fsm___pip_5160_1_94 = 0;
end
if ( (_ready_fsm___pip_5160_1_94)   && (_d__full_fsm___pip_5160_1_93)   && (!_t__stall_fsm___pip_5160_1_93)   && (!_d__full_fsm___pip_5160_1_94)   && (!_t__stall_fsm___pip_5160_1_94)   ) begin
   _d__idx_fsm___pip_5160_1_94 = 1;
   _d__full_fsm___pip_5160_1_93 = 0;
end
if ( (_ready_fsm___pip_5160_1_93)   && (_d__full_fsm___pip_5160_1_92)   && (!_t__stall_fsm___pip_5160_1_92)   && (!_d__full_fsm___pip_5160_1_93)   && (!_t__stall_fsm___pip_5160_1_93)   ) begin
   _d__idx_fsm___pip_5160_1_93 = 1;
   _d__full_fsm___pip_5160_1_92 = 0;
end
if ( (_ready_fsm___pip_5160_1_92)   && (_d__full_fsm___pip_5160_1_91)   && (!_t__stall_fsm___pip_5160_1_91)   && (!_d__full_fsm___pip_5160_1_92)   && (!_t__stall_fsm___pip_5160_1_92)   ) begin
   _d__idx_fsm___pip_5160_1_92 = 1;
   _d__full_fsm___pip_5160_1_91 = 0;
end
if ( (_ready_fsm___pip_5160_1_91)   && (_d__full_fsm___pip_5160_1_90)   && (!_t__stall_fsm___pip_5160_1_90)   && (!_d__full_fsm___pip_5160_1_91)   && (!_t__stall_fsm___pip_5160_1_91)   ) begin
   _d__idx_fsm___pip_5160_1_91 = 1;
   _d__full_fsm___pip_5160_1_90 = 0;
end
if ( (_ready_fsm___pip_5160_1_90)   && (_d__full_fsm___pip_5160_1_89)   && (!_t__stall_fsm___pip_5160_1_89)   && (!_d__full_fsm___pip_5160_1_90)   && (!_t__stall_fsm___pip_5160_1_90)   ) begin
   _d__idx_fsm___pip_5160_1_90 = 1;
   _d__full_fsm___pip_5160_1_89 = 0;
end
if ( (_ready_fsm___pip_5160_1_89)   && (_d__full_fsm___pip_5160_1_88)   && (!_t__stall_fsm___pip_5160_1_88)   && (!_d__full_fsm___pip_5160_1_89)   && (!_t__stall_fsm___pip_5160_1_89)   ) begin
   _d__idx_fsm___pip_5160_1_89 = 1;
   _d__full_fsm___pip_5160_1_88 = 0;
end
if ( (_ready_fsm___pip_5160_1_88)   && (_d__full_fsm___pip_5160_1_87)   && (!_t__stall_fsm___pip_5160_1_87)   && (!_d__full_fsm___pip_5160_1_88)   && (!_t__stall_fsm___pip_5160_1_88)   ) begin
   _d__idx_fsm___pip_5160_1_88 = 1;
   _d__full_fsm___pip_5160_1_87 = 0;
end
if ( (_ready_fsm___pip_5160_1_87)   && (_d__full_fsm___pip_5160_1_86)   && (!_t__stall_fsm___pip_5160_1_86)   && (!_d__full_fsm___pip_5160_1_87)   && (!_t__stall_fsm___pip_5160_1_87)   ) begin
   _d__idx_fsm___pip_5160_1_87 = 1;
   _d__full_fsm___pip_5160_1_86 = 0;
end
if ( (_ready_fsm___pip_5160_1_86)   && (_d__full_fsm___pip_5160_1_85)   && (!_t__stall_fsm___pip_5160_1_85)   && (!_d__full_fsm___pip_5160_1_86)   && (!_t__stall_fsm___pip_5160_1_86)   ) begin
   _d__idx_fsm___pip_5160_1_86 = 1;
   _d__full_fsm___pip_5160_1_85 = 0;
end
if ( (_ready_fsm___pip_5160_1_85)   && (_d__full_fsm___pip_5160_1_84)   && (!_t__stall_fsm___pip_5160_1_84)   && (!_d__full_fsm___pip_5160_1_85)   && (!_t__stall_fsm___pip_5160_1_85)   ) begin
   _d__idx_fsm___pip_5160_1_85 = 1;
   _d__full_fsm___pip_5160_1_84 = 0;
end
if ( (_ready_fsm___pip_5160_1_84)   && (_d__full_fsm___pip_5160_1_83)   && (!_t__stall_fsm___pip_5160_1_83)   && (!_d__full_fsm___pip_5160_1_84)   && (!_t__stall_fsm___pip_5160_1_84)   ) begin
   _d__idx_fsm___pip_5160_1_84 = 1;
   _d__full_fsm___pip_5160_1_83 = 0;
end
if ( (_ready_fsm___pip_5160_1_83)   && (_d__full_fsm___pip_5160_1_82)   && (!_t__stall_fsm___pip_5160_1_82)   && (!_d__full_fsm___pip_5160_1_83)   && (!_t__stall_fsm___pip_5160_1_83)   ) begin
   _d__idx_fsm___pip_5160_1_83 = 1;
   _d__full_fsm___pip_5160_1_82 = 0;
end
if ( (_ready_fsm___pip_5160_1_82)   && (_d__full_fsm___pip_5160_1_81)   && (!_t__stall_fsm___pip_5160_1_81)   && (!_d__full_fsm___pip_5160_1_82)   && (!_t__stall_fsm___pip_5160_1_82)   ) begin
   _d__idx_fsm___pip_5160_1_82 = 1;
   _d__full_fsm___pip_5160_1_81 = 0;
end
if ( (_ready_fsm___pip_5160_1_81)   && (_d__full_fsm___pip_5160_1_80)   && (!_t__stall_fsm___pip_5160_1_80)   && (!_d__full_fsm___pip_5160_1_81)   && (!_t__stall_fsm___pip_5160_1_81)   ) begin
   _d__idx_fsm___pip_5160_1_81 = 1;
   _d__full_fsm___pip_5160_1_80 = 0;
end
if ( (_ready_fsm___pip_5160_1_80)   && (_d__full_fsm___pip_5160_1_79)   && (!_t__stall_fsm___pip_5160_1_79)   && (!_d__full_fsm___pip_5160_1_80)   && (!_t__stall_fsm___pip_5160_1_80)   ) begin
   _d__idx_fsm___pip_5160_1_80 = 1;
   _d__full_fsm___pip_5160_1_79 = 0;
end
if ( (_ready_fsm___pip_5160_1_79)   && (_d__full_fsm___pip_5160_1_78)   && (!_t__stall_fsm___pip_5160_1_78)   && (!_d__full_fsm___pip_5160_1_79)   && (!_t__stall_fsm___pip_5160_1_79)   ) begin
   _d__idx_fsm___pip_5160_1_79 = 1;
   _d__full_fsm___pip_5160_1_78 = 0;
end
if ( (_ready_fsm___pip_5160_1_78)   && (_d__full_fsm___pip_5160_1_77)   && (!_t__stall_fsm___pip_5160_1_77)   && (!_d__full_fsm___pip_5160_1_78)   && (!_t__stall_fsm___pip_5160_1_78)   ) begin
   _d__idx_fsm___pip_5160_1_78 = 1;
   _d__full_fsm___pip_5160_1_77 = 0;
end
if ( (_ready_fsm___pip_5160_1_77)   && (_d__full_fsm___pip_5160_1_76)   && (!_t__stall_fsm___pip_5160_1_76)   && (!_d__full_fsm___pip_5160_1_77)   && (!_t__stall_fsm___pip_5160_1_77)   ) begin
   _d__idx_fsm___pip_5160_1_77 = 1;
   _d__full_fsm___pip_5160_1_76 = 0;
end
if ( (_ready_fsm___pip_5160_1_76)   && (_d__full_fsm___pip_5160_1_75)   && (!_t__stall_fsm___pip_5160_1_75)   && (!_d__full_fsm___pip_5160_1_76)   && (!_t__stall_fsm___pip_5160_1_76)   ) begin
   _d__idx_fsm___pip_5160_1_76 = 1;
   _d__full_fsm___pip_5160_1_75 = 0;
end
if ( (_ready_fsm___pip_5160_1_75)   && (_d__full_fsm___pip_5160_1_74)   && (!_t__stall_fsm___pip_5160_1_74)   && (!_d__full_fsm___pip_5160_1_75)   && (!_t__stall_fsm___pip_5160_1_75)   ) begin
   _d__idx_fsm___pip_5160_1_75 = 1;
   _d__full_fsm___pip_5160_1_74 = 0;
end
if ( (_ready_fsm___pip_5160_1_74)   && (_d__full_fsm___pip_5160_1_73)   && (!_t__stall_fsm___pip_5160_1_73)   && (!_d__full_fsm___pip_5160_1_74)   && (!_t__stall_fsm___pip_5160_1_74)   ) begin
   _d__idx_fsm___pip_5160_1_74 = 1;
   _d__full_fsm___pip_5160_1_73 = 0;
end
if ( (_ready_fsm___pip_5160_1_73)   && (_d__full_fsm___pip_5160_1_72)   && (!_t__stall_fsm___pip_5160_1_72)   && (!_d__full_fsm___pip_5160_1_73)   && (!_t__stall_fsm___pip_5160_1_73)   ) begin
   _d__idx_fsm___pip_5160_1_73 = 1;
   _d__full_fsm___pip_5160_1_72 = 0;
end
if ( (_ready_fsm___pip_5160_1_72)   && (_d__full_fsm___pip_5160_1_71)   && (!_t__stall_fsm___pip_5160_1_71)   && (!_d__full_fsm___pip_5160_1_72)   && (!_t__stall_fsm___pip_5160_1_72)   ) begin
   _d__idx_fsm___pip_5160_1_72 = 1;
   _d__full_fsm___pip_5160_1_71 = 0;
end
if ( (_ready_fsm___pip_5160_1_71)   && (_d__full_fsm___pip_5160_1_70)   && (!_t__stall_fsm___pip_5160_1_70)   && (!_d__full_fsm___pip_5160_1_71)   && (!_t__stall_fsm___pip_5160_1_71)   ) begin
   _d__idx_fsm___pip_5160_1_71 = 1;
   _d__full_fsm___pip_5160_1_70 = 0;
end
if ( (_ready_fsm___pip_5160_1_70)   && (_d__full_fsm___pip_5160_1_69)   && (!_t__stall_fsm___pip_5160_1_69)   && (!_d__full_fsm___pip_5160_1_70)   && (!_t__stall_fsm___pip_5160_1_70)   ) begin
   _d__idx_fsm___pip_5160_1_70 = 1;
   _d__full_fsm___pip_5160_1_69 = 0;
end
if ( (_ready_fsm___pip_5160_1_69)   && (_d__full_fsm___pip_5160_1_68)   && (!_t__stall_fsm___pip_5160_1_68)   && (!_d__full_fsm___pip_5160_1_69)   && (!_t__stall_fsm___pip_5160_1_69)   ) begin
   _d__idx_fsm___pip_5160_1_69 = 1;
   _d__full_fsm___pip_5160_1_68 = 0;
end
if ( (_ready_fsm___pip_5160_1_68)   && (_d__full_fsm___pip_5160_1_67)   && (!_t__stall_fsm___pip_5160_1_67)   && (!_d__full_fsm___pip_5160_1_68)   && (!_t__stall_fsm___pip_5160_1_68)   ) begin
   _d__idx_fsm___pip_5160_1_68 = 1;
   _d__full_fsm___pip_5160_1_67 = 0;
end
if ( (_ready_fsm___pip_5160_1_67)   && (_d__full_fsm___pip_5160_1_66)   && (!_t__stall_fsm___pip_5160_1_66)   && (!_d__full_fsm___pip_5160_1_67)   && (!_t__stall_fsm___pip_5160_1_67)   ) begin
   _d__idx_fsm___pip_5160_1_67 = 1;
   _d__full_fsm___pip_5160_1_66 = 0;
end
if ( (_ready_fsm___pip_5160_1_66)   && (_d__full_fsm___pip_5160_1_65)   && (!_t__stall_fsm___pip_5160_1_65)   && (!_d__full_fsm___pip_5160_1_66)   && (!_t__stall_fsm___pip_5160_1_66)   ) begin
   _d__idx_fsm___pip_5160_1_66 = 1;
   _d__full_fsm___pip_5160_1_65 = 0;
end
if ( (_ready_fsm___pip_5160_1_65)   && (_d__full_fsm___pip_5160_1_64)   && (!_t__stall_fsm___pip_5160_1_64)   && (!_d__full_fsm___pip_5160_1_65)   && (!_t__stall_fsm___pip_5160_1_65)   ) begin
   _d__idx_fsm___pip_5160_1_65 = 1;
   _d__full_fsm___pip_5160_1_64 = 0;
end
if ( (_ready_fsm___pip_5160_1_64)   && (_d__full_fsm___pip_5160_1_63)   && (!_t__stall_fsm___pip_5160_1_63)   && (!_d__full_fsm___pip_5160_1_64)   && (!_t__stall_fsm___pip_5160_1_64)   ) begin
   _d__idx_fsm___pip_5160_1_64 = 1;
   _d__full_fsm___pip_5160_1_63 = 0;
end
if ( (_ready_fsm___pip_5160_1_63)   && (_d__full_fsm___pip_5160_1_62)   && (!_t__stall_fsm___pip_5160_1_62)   && (!_d__full_fsm___pip_5160_1_63)   && (!_t__stall_fsm___pip_5160_1_63)   ) begin
   _d__idx_fsm___pip_5160_1_63 = 1;
   _d__full_fsm___pip_5160_1_62 = 0;
end
if ( (_ready_fsm___pip_5160_1_62)   && (_d__full_fsm___pip_5160_1_61)   && (!_t__stall_fsm___pip_5160_1_61)   && (!_d__full_fsm___pip_5160_1_62)   && (!_t__stall_fsm___pip_5160_1_62)   ) begin
   _d__idx_fsm___pip_5160_1_62 = 1;
   _d__full_fsm___pip_5160_1_61 = 0;
end
if ( (_ready_fsm___pip_5160_1_61)   && (_d__full_fsm___pip_5160_1_60)   && (!_t__stall_fsm___pip_5160_1_60)   && (!_d__full_fsm___pip_5160_1_61)   && (!_t__stall_fsm___pip_5160_1_61)   ) begin
   _d__idx_fsm___pip_5160_1_61 = 1;
   _d__full_fsm___pip_5160_1_60 = 0;
end
if ( (_ready_fsm___pip_5160_1_60)   && (_d__full_fsm___pip_5160_1_59)   && (!_t__stall_fsm___pip_5160_1_59)   && (!_d__full_fsm___pip_5160_1_60)   && (!_t__stall_fsm___pip_5160_1_60)   ) begin
   _d__idx_fsm___pip_5160_1_60 = 1;
   _d__full_fsm___pip_5160_1_59 = 0;
end
if ( (_ready_fsm___pip_5160_1_59)   && (_d__full_fsm___pip_5160_1_58)   && (!_t__stall_fsm___pip_5160_1_58)   && (!_d__full_fsm___pip_5160_1_59)   && (!_t__stall_fsm___pip_5160_1_59)   ) begin
   _d__idx_fsm___pip_5160_1_59 = 1;
   _d__full_fsm___pip_5160_1_58 = 0;
end
if ( (_ready_fsm___pip_5160_1_58)   && (_d__full_fsm___pip_5160_1_57)   && (!_t__stall_fsm___pip_5160_1_57)   && (!_d__full_fsm___pip_5160_1_58)   && (!_t__stall_fsm___pip_5160_1_58)   ) begin
   _d__idx_fsm___pip_5160_1_58 = 1;
   _d__full_fsm___pip_5160_1_57 = 0;
end
if ( (_ready_fsm___pip_5160_1_57)   && (_d__full_fsm___pip_5160_1_56)   && (!_t__stall_fsm___pip_5160_1_56)   && (!_d__full_fsm___pip_5160_1_57)   && (!_t__stall_fsm___pip_5160_1_57)   ) begin
   _d__idx_fsm___pip_5160_1_57 = 1;
   _d__full_fsm___pip_5160_1_56 = 0;
end
if ( (_ready_fsm___pip_5160_1_56)   && (_d__full_fsm___pip_5160_1_55)   && (!_t__stall_fsm___pip_5160_1_55)   && (!_d__full_fsm___pip_5160_1_56)   && (!_t__stall_fsm___pip_5160_1_56)   ) begin
   _d__idx_fsm___pip_5160_1_56 = 1;
   _d__full_fsm___pip_5160_1_55 = 0;
end
if ( (_ready_fsm___pip_5160_1_55)   && (_d__full_fsm___pip_5160_1_54)   && (!_t__stall_fsm___pip_5160_1_54)   && (!_d__full_fsm___pip_5160_1_55)   && (!_t__stall_fsm___pip_5160_1_55)   ) begin
   _d__idx_fsm___pip_5160_1_55 = 1;
   _d__full_fsm___pip_5160_1_54 = 0;
end
if ( (_ready_fsm___pip_5160_1_54)   && (_d__full_fsm___pip_5160_1_53)   && (!_t__stall_fsm___pip_5160_1_53)   && (!_d__full_fsm___pip_5160_1_54)   && (!_t__stall_fsm___pip_5160_1_54)   ) begin
   _d__idx_fsm___pip_5160_1_54 = 1;
   _d__full_fsm___pip_5160_1_53 = 0;
end
if ( (_ready_fsm___pip_5160_1_53)   && (_d__full_fsm___pip_5160_1_52)   && (!_t__stall_fsm___pip_5160_1_52)   && (!_d__full_fsm___pip_5160_1_53)   && (!_t__stall_fsm___pip_5160_1_53)   ) begin
   _d__idx_fsm___pip_5160_1_53 = 1;
   _d__full_fsm___pip_5160_1_52 = 0;
end
if ( (_ready_fsm___pip_5160_1_52)   && (_d__full_fsm___pip_5160_1_51)   && (!_t__stall_fsm___pip_5160_1_51)   && (!_d__full_fsm___pip_5160_1_52)   && (!_t__stall_fsm___pip_5160_1_52)   ) begin
   _d__idx_fsm___pip_5160_1_52 = 1;
   _d__full_fsm___pip_5160_1_51 = 0;
end
if ( (_ready_fsm___pip_5160_1_51)   && (_d__full_fsm___pip_5160_1_50)   && (!_t__stall_fsm___pip_5160_1_50)   && (!_d__full_fsm___pip_5160_1_51)   && (!_t__stall_fsm___pip_5160_1_51)   ) begin
   _d__idx_fsm___pip_5160_1_51 = 1;
   _d__full_fsm___pip_5160_1_50 = 0;
end
if ( (_ready_fsm___pip_5160_1_50)   && (_d__full_fsm___pip_5160_1_49)   && (!_t__stall_fsm___pip_5160_1_49)   && (!_d__full_fsm___pip_5160_1_50)   && (!_t__stall_fsm___pip_5160_1_50)   ) begin
   _d__idx_fsm___pip_5160_1_50 = 1;
   _d__full_fsm___pip_5160_1_49 = 0;
end
if ( (_ready_fsm___pip_5160_1_49)   && (_d__full_fsm___pip_5160_1_48)   && (!_t__stall_fsm___pip_5160_1_48)   && (!_d__full_fsm___pip_5160_1_49)   && (!_t__stall_fsm___pip_5160_1_49)   ) begin
   _d__idx_fsm___pip_5160_1_49 = 1;
   _d__full_fsm___pip_5160_1_48 = 0;
end
if ( (_ready_fsm___pip_5160_1_48)   && (_d__full_fsm___pip_5160_1_47)   && (!_t__stall_fsm___pip_5160_1_47)   && (!_d__full_fsm___pip_5160_1_48)   && (!_t__stall_fsm___pip_5160_1_48)   ) begin
   _d__idx_fsm___pip_5160_1_48 = 1;
   _d__full_fsm___pip_5160_1_47 = 0;
end
if ( (_ready_fsm___pip_5160_1_47)   && (_d__full_fsm___pip_5160_1_46)   && (!_t__stall_fsm___pip_5160_1_46)   && (!_d__full_fsm___pip_5160_1_47)   && (!_t__stall_fsm___pip_5160_1_47)   ) begin
   _d__idx_fsm___pip_5160_1_47 = 1;
   _d__full_fsm___pip_5160_1_46 = 0;
end
if ( (_ready_fsm___pip_5160_1_46)   && (_d__full_fsm___pip_5160_1_45)   && (!_t__stall_fsm___pip_5160_1_45)   && (!_d__full_fsm___pip_5160_1_46)   && (!_t__stall_fsm___pip_5160_1_46)   ) begin
   _d__idx_fsm___pip_5160_1_46 = 1;
   _d__full_fsm___pip_5160_1_45 = 0;
end
if ( (_ready_fsm___pip_5160_1_45)   && (_d__full_fsm___pip_5160_1_44)   && (!_t__stall_fsm___pip_5160_1_44)   && (!_d__full_fsm___pip_5160_1_45)   && (!_t__stall_fsm___pip_5160_1_45)   ) begin
   _d__idx_fsm___pip_5160_1_45 = 1;
   _d__full_fsm___pip_5160_1_44 = 0;
end
if ( (_ready_fsm___pip_5160_1_44)   && (_d__full_fsm___pip_5160_1_43)   && (!_t__stall_fsm___pip_5160_1_43)   && (!_d__full_fsm___pip_5160_1_44)   && (!_t__stall_fsm___pip_5160_1_44)   ) begin
   _d__idx_fsm___pip_5160_1_44 = 1;
   _d__full_fsm___pip_5160_1_43 = 0;
end
if ( (_ready_fsm___pip_5160_1_43)   && (_d__full_fsm___pip_5160_1_42)   && (!_t__stall_fsm___pip_5160_1_42)   && (!_d__full_fsm___pip_5160_1_43)   && (!_t__stall_fsm___pip_5160_1_43)   ) begin
   _d__idx_fsm___pip_5160_1_43 = 1;
   _d__full_fsm___pip_5160_1_42 = 0;
end
if ( (_ready_fsm___pip_5160_1_42)   && (_d__full_fsm___pip_5160_1_41)   && (!_t__stall_fsm___pip_5160_1_41)   && (!_d__full_fsm___pip_5160_1_42)   && (!_t__stall_fsm___pip_5160_1_42)   ) begin
   _d__idx_fsm___pip_5160_1_42 = 1;
   _d__full_fsm___pip_5160_1_41 = 0;
end
if ( (_ready_fsm___pip_5160_1_41)   && (_d__full_fsm___pip_5160_1_40)   && (!_t__stall_fsm___pip_5160_1_40)   && (!_d__full_fsm___pip_5160_1_41)   && (!_t__stall_fsm___pip_5160_1_41)   ) begin
   _d__idx_fsm___pip_5160_1_41 = 1;
   _d__full_fsm___pip_5160_1_40 = 0;
end
if ( (_ready_fsm___pip_5160_1_40)   && (_d__full_fsm___pip_5160_1_39)   && (!_t__stall_fsm___pip_5160_1_39)   && (!_d__full_fsm___pip_5160_1_40)   && (!_t__stall_fsm___pip_5160_1_40)   ) begin
   _d__idx_fsm___pip_5160_1_40 = 1;
   _d__full_fsm___pip_5160_1_39 = 0;
end
if ( (_ready_fsm___pip_5160_1_39)   && (_d__full_fsm___pip_5160_1_38)   && (!_t__stall_fsm___pip_5160_1_38)   && (!_d__full_fsm___pip_5160_1_39)   && (!_t__stall_fsm___pip_5160_1_39)   ) begin
   _d__idx_fsm___pip_5160_1_39 = 1;
   _d__full_fsm___pip_5160_1_38 = 0;
end
if ( (_ready_fsm___pip_5160_1_38)   && (_d__full_fsm___pip_5160_1_37)   && (!_t__stall_fsm___pip_5160_1_37)   && (!_d__full_fsm___pip_5160_1_38)   && (!_t__stall_fsm___pip_5160_1_38)   ) begin
   _d__idx_fsm___pip_5160_1_38 = 1;
   _d__full_fsm___pip_5160_1_37 = 0;
end
if ( (_ready_fsm___pip_5160_1_37)   && (_d__full_fsm___pip_5160_1_36)   && (!_t__stall_fsm___pip_5160_1_36)   && (!_d__full_fsm___pip_5160_1_37)   && (!_t__stall_fsm___pip_5160_1_37)   ) begin
   _d__idx_fsm___pip_5160_1_37 = 1;
   _d__full_fsm___pip_5160_1_36 = 0;
end
if ( (_ready_fsm___pip_5160_1_36)   && (_d__full_fsm___pip_5160_1_35)   && (!_t__stall_fsm___pip_5160_1_35)   && (!_d__full_fsm___pip_5160_1_36)   && (!_t__stall_fsm___pip_5160_1_36)   ) begin
   _d__idx_fsm___pip_5160_1_36 = 1;
   _d__full_fsm___pip_5160_1_35 = 0;
end
if ( (_ready_fsm___pip_5160_1_35)   && (_d__full_fsm___pip_5160_1_34)   && (!_t__stall_fsm___pip_5160_1_34)   && (!_d__full_fsm___pip_5160_1_35)   && (!_t__stall_fsm___pip_5160_1_35)   ) begin
   _d__idx_fsm___pip_5160_1_35 = 1;
   _d__full_fsm___pip_5160_1_34 = 0;
end
if ( (_ready_fsm___pip_5160_1_34)   && (_d__full_fsm___pip_5160_1_33)   && (!_t__stall_fsm___pip_5160_1_33)   && (!_d__full_fsm___pip_5160_1_34)   && (!_t__stall_fsm___pip_5160_1_34)   ) begin
   _d__idx_fsm___pip_5160_1_34 = 1;
   _d__full_fsm___pip_5160_1_33 = 0;
end
if ( (_ready_fsm___pip_5160_1_33)   && (_d__full_fsm___pip_5160_1_32)   && (!_t__stall_fsm___pip_5160_1_32)   && (!_d__full_fsm___pip_5160_1_33)   && (!_t__stall_fsm___pip_5160_1_33)   ) begin
   _d__idx_fsm___pip_5160_1_33 = 1;
   _d__full_fsm___pip_5160_1_32 = 0;
end
if ( (_ready_fsm___pip_5160_1_32)   && (_d__full_fsm___pip_5160_1_31)   && (!_t__stall_fsm___pip_5160_1_31)   && (!_d__full_fsm___pip_5160_1_32)   && (!_t__stall_fsm___pip_5160_1_32)   ) begin
   _d__idx_fsm___pip_5160_1_32 = 1;
   _d__full_fsm___pip_5160_1_31 = 0;
end
if ( (_ready_fsm___pip_5160_1_31)   && (_d__full_fsm___pip_5160_1_30)   && (!_t__stall_fsm___pip_5160_1_30)   && (!_d__full_fsm___pip_5160_1_31)   && (!_t__stall_fsm___pip_5160_1_31)   ) begin
   _d__idx_fsm___pip_5160_1_31 = 1;
   _d__full_fsm___pip_5160_1_30 = 0;
end
if ( (_ready_fsm___pip_5160_1_30)   && (_d__full_fsm___pip_5160_1_29)   && (!_t__stall_fsm___pip_5160_1_29)   && (!_d__full_fsm___pip_5160_1_30)   && (!_t__stall_fsm___pip_5160_1_30)   ) begin
   _d__idx_fsm___pip_5160_1_30 = 1;
   _d__full_fsm___pip_5160_1_29 = 0;
end
if ( (_ready_fsm___pip_5160_1_29)   && (_d__full_fsm___pip_5160_1_28)   && (!_t__stall_fsm___pip_5160_1_28)   && (!_d__full_fsm___pip_5160_1_29)   && (!_t__stall_fsm___pip_5160_1_29)   ) begin
   _d__idx_fsm___pip_5160_1_29 = 1;
   _d__full_fsm___pip_5160_1_28 = 0;
end
if ( (_ready_fsm___pip_5160_1_28)   && (_d__full_fsm___pip_5160_1_27)   && (!_t__stall_fsm___pip_5160_1_27)   && (!_d__full_fsm___pip_5160_1_28)   && (!_t__stall_fsm___pip_5160_1_28)   ) begin
   _d__idx_fsm___pip_5160_1_28 = 1;
   _d__full_fsm___pip_5160_1_27 = 0;
end
if ( (_ready_fsm___pip_5160_1_27)   && (_d__full_fsm___pip_5160_1_26)   && (!_t__stall_fsm___pip_5160_1_26)   && (!_d__full_fsm___pip_5160_1_27)   && (!_t__stall_fsm___pip_5160_1_27)   ) begin
   _d__idx_fsm___pip_5160_1_27 = 1;
   _d__full_fsm___pip_5160_1_26 = 0;
end
if ( (_ready_fsm___pip_5160_1_26)   && (_d__full_fsm___pip_5160_1_25)   && (!_t__stall_fsm___pip_5160_1_25)   && (!_d__full_fsm___pip_5160_1_26)   && (!_t__stall_fsm___pip_5160_1_26)   ) begin
   _d__idx_fsm___pip_5160_1_26 = 1;
   _d__full_fsm___pip_5160_1_25 = 0;
end
if ( (_ready_fsm___pip_5160_1_25)   && (_d__full_fsm___pip_5160_1_24)   && (!_t__stall_fsm___pip_5160_1_24)   && (!_d__full_fsm___pip_5160_1_25)   && (!_t__stall_fsm___pip_5160_1_25)   ) begin
   _d__idx_fsm___pip_5160_1_25 = 1;
   _d__full_fsm___pip_5160_1_24 = 0;
end
if ( (_ready_fsm___pip_5160_1_24)   && (_d__full_fsm___pip_5160_1_23)   && (!_t__stall_fsm___pip_5160_1_23)   && (!_d__full_fsm___pip_5160_1_24)   && (!_t__stall_fsm___pip_5160_1_24)   ) begin
   _d__idx_fsm___pip_5160_1_24 = 1;
   _d__full_fsm___pip_5160_1_23 = 0;
end
if ( (_ready_fsm___pip_5160_1_23)   && (_d__full_fsm___pip_5160_1_22)   && (!_t__stall_fsm___pip_5160_1_22)   && (!_d__full_fsm___pip_5160_1_23)   && (!_t__stall_fsm___pip_5160_1_23)   ) begin
   _d__idx_fsm___pip_5160_1_23 = 1;
   _d__full_fsm___pip_5160_1_22 = 0;
end
if ( (_ready_fsm___pip_5160_1_22)   && (_d__full_fsm___pip_5160_1_21)   && (!_t__stall_fsm___pip_5160_1_21)   && (!_d__full_fsm___pip_5160_1_22)   && (!_t__stall_fsm___pip_5160_1_22)   ) begin
   _d__idx_fsm___pip_5160_1_22 = 1;
   _d__full_fsm___pip_5160_1_21 = 0;
end
if ( (_ready_fsm___pip_5160_1_21)   && (_d__full_fsm___pip_5160_1_20)   && (!_t__stall_fsm___pip_5160_1_20)   && (!_d__full_fsm___pip_5160_1_21)   && (!_t__stall_fsm___pip_5160_1_21)   ) begin
   _d__idx_fsm___pip_5160_1_21 = 1;
   _d__full_fsm___pip_5160_1_20 = 0;
end
if ( (_ready_fsm___pip_5160_1_20)   && (_d__full_fsm___pip_5160_1_19)   && (!_t__stall_fsm___pip_5160_1_19)   && (!_d__full_fsm___pip_5160_1_20)   && (!_t__stall_fsm___pip_5160_1_20)   ) begin
   _d__idx_fsm___pip_5160_1_20 = 1;
   _d__full_fsm___pip_5160_1_19 = 0;
end
if ( (_ready_fsm___pip_5160_1_19)   && (_d__full_fsm___pip_5160_1_18)   && (!_t__stall_fsm___pip_5160_1_18)   && (!_d__full_fsm___pip_5160_1_19)   && (!_t__stall_fsm___pip_5160_1_19)   ) begin
   _d__idx_fsm___pip_5160_1_19 = 1;
   _d__full_fsm___pip_5160_1_18 = 0;
end
if ( (_ready_fsm___pip_5160_1_18)   && (_d__full_fsm___pip_5160_1_17)   && (!_t__stall_fsm___pip_5160_1_17)   && (!_d__full_fsm___pip_5160_1_18)   && (!_t__stall_fsm___pip_5160_1_18)   ) begin
   _d__idx_fsm___pip_5160_1_18 = 1;
   _d__full_fsm___pip_5160_1_17 = 0;
end
if ( (_ready_fsm___pip_5160_1_17)   && (_d__full_fsm___pip_5160_1_16)   && (!_t__stall_fsm___pip_5160_1_16)   && (!_d__full_fsm___pip_5160_1_17)   && (!_t__stall_fsm___pip_5160_1_17)   ) begin
   _d__idx_fsm___pip_5160_1_17 = 1;
   _d__full_fsm___pip_5160_1_16 = 0;
end
if ( (_ready_fsm___pip_5160_1_16)   && (_d__full_fsm___pip_5160_1_15)   && (!_t__stall_fsm___pip_5160_1_15)   && (!_d__full_fsm___pip_5160_1_16)   && (!_t__stall_fsm___pip_5160_1_16)   ) begin
   _d__idx_fsm___pip_5160_1_16 = 1;
   _d__full_fsm___pip_5160_1_15 = 0;
end
if ( (_ready_fsm___pip_5160_1_15)   && (_d__full_fsm___pip_5160_1_14)   && (!_t__stall_fsm___pip_5160_1_14)   && (!_d__full_fsm___pip_5160_1_15)   && (!_t__stall_fsm___pip_5160_1_15)   ) begin
   _d__idx_fsm___pip_5160_1_15 = 1;
   _d__full_fsm___pip_5160_1_14 = 0;
end
if ( (_ready_fsm___pip_5160_1_14)   && (_d__full_fsm___pip_5160_1_13)   && (!_t__stall_fsm___pip_5160_1_13)   && (!_d__full_fsm___pip_5160_1_14)   && (!_t__stall_fsm___pip_5160_1_14)   ) begin
   _d__idx_fsm___pip_5160_1_14 = 1;
   _d__full_fsm___pip_5160_1_13 = 0;
end
if ( (_ready_fsm___pip_5160_1_13)   && (_d__full_fsm___pip_5160_1_12)   && (!_t__stall_fsm___pip_5160_1_12)   && (!_d__full_fsm___pip_5160_1_13)   && (!_t__stall_fsm___pip_5160_1_13)   ) begin
   _d__idx_fsm___pip_5160_1_13 = 1;
   _d__full_fsm___pip_5160_1_12 = 0;
end
if ( (_ready_fsm___pip_5160_1_12)   && (_d__full_fsm___pip_5160_1_11)   && (!_t__stall_fsm___pip_5160_1_11)   && (!_d__full_fsm___pip_5160_1_12)   && (!_t__stall_fsm___pip_5160_1_12)   ) begin
   _d__idx_fsm___pip_5160_1_12 = 1;
   _d__full_fsm___pip_5160_1_11 = 0;
end
if ( (_ready_fsm___pip_5160_1_11)   && (_d__full_fsm___pip_5160_1_10)   && (!_t__stall_fsm___pip_5160_1_10)   && (!_d__full_fsm___pip_5160_1_11)   && (!_t__stall_fsm___pip_5160_1_11)   ) begin
   _d__idx_fsm___pip_5160_1_11 = 1;
   _d__full_fsm___pip_5160_1_10 = 0;
end
if ( (_ready_fsm___pip_5160_1_10)   && (_d__full_fsm___pip_5160_1_9)   && (!_t__stall_fsm___pip_5160_1_9)   && (!_d__full_fsm___pip_5160_1_10)   && (!_t__stall_fsm___pip_5160_1_10)   ) begin
   _d__idx_fsm___pip_5160_1_10 = 1;
   _d__full_fsm___pip_5160_1_9 = 0;
end
if ( (_ready_fsm___pip_5160_1_9)   && (_d__full_fsm___pip_5160_1_8)   && (!_t__stall_fsm___pip_5160_1_8)   && (!_d__full_fsm___pip_5160_1_9)   && (!_t__stall_fsm___pip_5160_1_9)   ) begin
   _d__idx_fsm___pip_5160_1_9 = 1;
   _d__full_fsm___pip_5160_1_8 = 0;
end
if ( (_ready_fsm___pip_5160_1_8)   && (_d__full_fsm___pip_5160_1_7)   && (!_t__stall_fsm___pip_5160_1_7)   && (!_d__full_fsm___pip_5160_1_8)   && (!_t__stall_fsm___pip_5160_1_8)   ) begin
   _d__idx_fsm___pip_5160_1_8 = 1;
   _d__full_fsm___pip_5160_1_7 = 0;
end
if ( (_ready_fsm___pip_5160_1_7)   && (_d__full_fsm___pip_5160_1_6)   && (!_t__stall_fsm___pip_5160_1_6)   && (!_d__full_fsm___pip_5160_1_7)   && (!_t__stall_fsm___pip_5160_1_7)   ) begin
   _d__idx_fsm___pip_5160_1_7 = 1;
   _d__full_fsm___pip_5160_1_6 = 0;
end
if ( (_ready_fsm___pip_5160_1_6)   && (_d__full_fsm___pip_5160_1_5)   && (!_t__stall_fsm___pip_5160_1_5)   && (!_d__full_fsm___pip_5160_1_6)   && (!_t__stall_fsm___pip_5160_1_6)   ) begin
   _d__idx_fsm___pip_5160_1_6 = 1;
   _d__full_fsm___pip_5160_1_5 = 0;
end
if ( (_ready_fsm___pip_5160_1_5)   && (_d__full_fsm___pip_5160_1_4)   && (!_t__stall_fsm___pip_5160_1_4)   && (!_d__full_fsm___pip_5160_1_5)   && (!_t__stall_fsm___pip_5160_1_5)   ) begin
   _d__idx_fsm___pip_5160_1_5 = 1;
   _d__full_fsm___pip_5160_1_4 = 0;
end
if ( (_ready_fsm___pip_5160_1_4)   && (_d__full_fsm___pip_5160_1_3)   && (!_t__stall_fsm___pip_5160_1_3)   && (!_d__full_fsm___pip_5160_1_4)   && (!_t__stall_fsm___pip_5160_1_4)   ) begin
   _d__idx_fsm___pip_5160_1_4 = 1;
   _d__full_fsm___pip_5160_1_3 = 0;
end
if ( (_ready_fsm___pip_5160_1_3)   && (_d__full_fsm___pip_5160_1_2)   && (!_t__stall_fsm___pip_5160_1_2)   && (!_d__full_fsm___pip_5160_1_3)   && (!_t__stall_fsm___pip_5160_1_3)   ) begin
   _d__idx_fsm___pip_5160_1_3 = 1;
   _d__full_fsm___pip_5160_1_2 = 0;
end
if ( (_ready_fsm___pip_5160_1_2)   && (_d__full_fsm___pip_5160_1_1)   && (!_t__stall_fsm___pip_5160_1_1)   && (!_d__full_fsm___pip_5160_1_2)   && (!_t__stall_fsm___pip_5160_1_2)   ) begin
   _d__idx_fsm___pip_5160_1_2 = 1;
   _d__full_fsm___pip_5160_1_1 = 0;
end
if ( (_ready_fsm___pip_5160_1_1)   && (_d__full_fsm___pip_5160_1_0)   && (!_t__stall_fsm___pip_5160_1_0)   && (!_d__full_fsm___pip_5160_1_1)   && (!_t__stall_fsm___pip_5160_1_1)   ) begin
   _d__idx_fsm___pip_5160_1_1 = 1;
   _d__full_fsm___pip_5160_1_0 = 0;
end
if ( (_ready_fsm___pip_5160_1_0)   && ((( ~_autorun ? 1 : _d__idx_fsm0)) == 2)
  && (!_d__full_fsm___pip_5160_1_0)   && (!_t__stall_fsm___pip_5160_1_0)   ) begin
   _d__idx_fsm___pip_5160_1_0 = 1;
end
end

always @(posedge clock) begin
_q_frame <= _d_frame;
_q_cos_addr0 <= _d_cos_addr0;
_q_cos_addr1 <= _d_cos_addr1;
_q_sin_addr0 <= _d_sin_addr0;
_q_sin_addr1 <= _d_sin_addr1;
_q_invA_addr0 <= _d_invA_addr0;
_q_invA_addr1 <= _d_invA_addr1;
_q_invB_addr <= _d_invB_addr;
_q___pip_5160_1_3___block_25_r_x_delta <= _d___pip_5160_1_3___block_25_r_x_delta;
_q___pip_5160_1_4___block_25_r_x_delta <= (_d__idx_fsm___pip_5160_1_4 == 1 && !_t__stall_fsm___pip_5160_1_4) ? _d___pip_5160_1_3___block_25_r_x_delta : _d___pip_5160_1_4___block_25_r_x_delta;
_q___pip_5160_1_3___block_25_r_z_delta <= _d___pip_5160_1_3___block_25_r_z_delta;
_q___pip_5160_1_4___block_25_r_z_delta <= (_d__idx_fsm___pip_5160_1_4 == 1 && !_t__stall_fsm___pip_5160_1_4) ? _d___pip_5160_1_3___block_25_r_z_delta : _d___pip_5160_1_4___block_25_r_z_delta;
_q___pip_5160_1_135___block_2731_clr_b <= _d___pip_5160_1_135___block_2731_clr_b;
_q___pip_5160_1_136___block_2731_clr_b <= (_d__idx_fsm___pip_5160_1_136 == 1 && !_t__stall_fsm___pip_5160_1_136) ? _d___pip_5160_1_135___block_2731_clr_b : _d___pip_5160_1_136___block_2731_clr_b;
_q___pip_5160_1_135___block_2731_clr_g <= _d___pip_5160_1_135___block_2731_clr_g;
_q___pip_5160_1_136___block_2731_clr_g <= (_d__idx_fsm___pip_5160_1_136 == 1 && !_t__stall_fsm___pip_5160_1_136) ? _d___pip_5160_1_135___block_2731_clr_g : _d___pip_5160_1_136___block_2731_clr_g;
_q___pip_5160_1_135___block_2731_clr_r <= _d___pip_5160_1_135___block_2731_clr_r;
_q___pip_5160_1_136___block_2731_clr_r <= (_d__idx_fsm___pip_5160_1_136 == 1 && !_t__stall_fsm___pip_5160_1_136) ? _d___pip_5160_1_135___block_2731_clr_r : _d___pip_5160_1_136___block_2731_clr_r;
_q___pip_5160_1_6___block_34_tm_x <= _d___pip_5160_1_6___block_34_tm_x;
_q___pip_5160_1_7___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___block_34_tm_x : _d___pip_5160_1_7___block_34_tm_x;
_q___pip_5160_1_8___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___block_34_tm_x : _d___pip_5160_1_8___block_34_tm_x;
_q___pip_5160_1_9___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___block_34_tm_x : _d___pip_5160_1_9___block_34_tm_x;
_q___pip_5160_1_10___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___block_34_tm_x : _d___pip_5160_1_10___block_34_tm_x;
_q___pip_5160_1_11___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___block_34_tm_x : _d___pip_5160_1_11___block_34_tm_x;
_q___pip_5160_1_12___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___block_34_tm_x : _d___pip_5160_1_12___block_34_tm_x;
_q___pip_5160_1_13___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___block_34_tm_x : _d___pip_5160_1_13___block_34_tm_x;
_q___pip_5160_1_14___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___block_34_tm_x : _d___pip_5160_1_14___block_34_tm_x;
_q___pip_5160_1_15___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___block_34_tm_x : _d___pip_5160_1_15___block_34_tm_x;
_q___pip_5160_1_16___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___block_34_tm_x : _d___pip_5160_1_16___block_34_tm_x;
_q___pip_5160_1_17___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___block_34_tm_x : _d___pip_5160_1_17___block_34_tm_x;
_q___pip_5160_1_18___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___block_34_tm_x : _d___pip_5160_1_18___block_34_tm_x;
_q___pip_5160_1_19___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___block_34_tm_x : _d___pip_5160_1_19___block_34_tm_x;
_q___pip_5160_1_20___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___block_34_tm_x : _d___pip_5160_1_20___block_34_tm_x;
_q___pip_5160_1_21___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___block_34_tm_x : _d___pip_5160_1_21___block_34_tm_x;
_q___pip_5160_1_22___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___block_34_tm_x : _d___pip_5160_1_22___block_34_tm_x;
_q___pip_5160_1_23___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___block_34_tm_x : _d___pip_5160_1_23___block_34_tm_x;
_q___pip_5160_1_24___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___block_34_tm_x : _d___pip_5160_1_24___block_34_tm_x;
_q___pip_5160_1_25___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___block_34_tm_x : _d___pip_5160_1_25___block_34_tm_x;
_q___pip_5160_1_26___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___block_34_tm_x : _d___pip_5160_1_26___block_34_tm_x;
_q___pip_5160_1_27___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___block_34_tm_x : _d___pip_5160_1_27___block_34_tm_x;
_q___pip_5160_1_28___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___block_34_tm_x : _d___pip_5160_1_28___block_34_tm_x;
_q___pip_5160_1_29___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___block_34_tm_x : _d___pip_5160_1_29___block_34_tm_x;
_q___pip_5160_1_30___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___block_34_tm_x : _d___pip_5160_1_30___block_34_tm_x;
_q___pip_5160_1_31___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___block_34_tm_x : _d___pip_5160_1_31___block_34_tm_x;
_q___pip_5160_1_32___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___block_34_tm_x : _d___pip_5160_1_32___block_34_tm_x;
_q___pip_5160_1_33___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___block_34_tm_x : _d___pip_5160_1_33___block_34_tm_x;
_q___pip_5160_1_34___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___block_34_tm_x : _d___pip_5160_1_34___block_34_tm_x;
_q___pip_5160_1_35___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___block_34_tm_x : _d___pip_5160_1_35___block_34_tm_x;
_q___pip_5160_1_36___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___block_34_tm_x : _d___pip_5160_1_36___block_34_tm_x;
_q___pip_5160_1_37___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___block_34_tm_x : _d___pip_5160_1_37___block_34_tm_x;
_q___pip_5160_1_38___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___block_34_tm_x : _d___pip_5160_1_38___block_34_tm_x;
_q___pip_5160_1_39___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___block_34_tm_x : _d___pip_5160_1_39___block_34_tm_x;
_q___pip_5160_1_40___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___block_34_tm_x : _d___pip_5160_1_40___block_34_tm_x;
_q___pip_5160_1_41___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___block_34_tm_x : _d___pip_5160_1_41___block_34_tm_x;
_q___pip_5160_1_42___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___block_34_tm_x : _d___pip_5160_1_42___block_34_tm_x;
_q___pip_5160_1_43___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___block_34_tm_x : _d___pip_5160_1_43___block_34_tm_x;
_q___pip_5160_1_44___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___block_34_tm_x : _d___pip_5160_1_44___block_34_tm_x;
_q___pip_5160_1_45___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___block_34_tm_x : _d___pip_5160_1_45___block_34_tm_x;
_q___pip_5160_1_46___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___block_34_tm_x : _d___pip_5160_1_46___block_34_tm_x;
_q___pip_5160_1_47___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___block_34_tm_x : _d___pip_5160_1_47___block_34_tm_x;
_q___pip_5160_1_48___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___block_34_tm_x : _d___pip_5160_1_48___block_34_tm_x;
_q___pip_5160_1_49___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___block_34_tm_x : _d___pip_5160_1_49___block_34_tm_x;
_q___pip_5160_1_50___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___block_34_tm_x : _d___pip_5160_1_50___block_34_tm_x;
_q___pip_5160_1_51___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___block_34_tm_x : _d___pip_5160_1_51___block_34_tm_x;
_q___pip_5160_1_52___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___block_34_tm_x : _d___pip_5160_1_52___block_34_tm_x;
_q___pip_5160_1_53___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___block_34_tm_x : _d___pip_5160_1_53___block_34_tm_x;
_q___pip_5160_1_54___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___block_34_tm_x : _d___pip_5160_1_54___block_34_tm_x;
_q___pip_5160_1_55___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___block_34_tm_x : _d___pip_5160_1_55___block_34_tm_x;
_q___pip_5160_1_56___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___block_34_tm_x : _d___pip_5160_1_56___block_34_tm_x;
_q___pip_5160_1_57___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___block_34_tm_x : _d___pip_5160_1_57___block_34_tm_x;
_q___pip_5160_1_58___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___block_34_tm_x : _d___pip_5160_1_58___block_34_tm_x;
_q___pip_5160_1_59___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___block_34_tm_x : _d___pip_5160_1_59___block_34_tm_x;
_q___pip_5160_1_60___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___block_34_tm_x : _d___pip_5160_1_60___block_34_tm_x;
_q___pip_5160_1_61___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___block_34_tm_x : _d___pip_5160_1_61___block_34_tm_x;
_q___pip_5160_1_62___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___block_34_tm_x : _d___pip_5160_1_62___block_34_tm_x;
_q___pip_5160_1_63___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___block_34_tm_x : _d___pip_5160_1_63___block_34_tm_x;
_q___pip_5160_1_64___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___block_34_tm_x : _d___pip_5160_1_64___block_34_tm_x;
_q___pip_5160_1_65___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___block_34_tm_x : _d___pip_5160_1_65___block_34_tm_x;
_q___pip_5160_1_66___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___block_34_tm_x : _d___pip_5160_1_66___block_34_tm_x;
_q___pip_5160_1_67___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___block_34_tm_x : _d___pip_5160_1_67___block_34_tm_x;
_q___pip_5160_1_68___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___block_34_tm_x : _d___pip_5160_1_68___block_34_tm_x;
_q___pip_5160_1_69___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___block_34_tm_x : _d___pip_5160_1_69___block_34_tm_x;
_q___pip_5160_1_70___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___block_34_tm_x : _d___pip_5160_1_70___block_34_tm_x;
_q___pip_5160_1_71___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___block_34_tm_x : _d___pip_5160_1_71___block_34_tm_x;
_q___pip_5160_1_72___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___block_34_tm_x : _d___pip_5160_1_72___block_34_tm_x;
_q___pip_5160_1_73___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___block_34_tm_x : _d___pip_5160_1_73___block_34_tm_x;
_q___pip_5160_1_74___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___block_34_tm_x : _d___pip_5160_1_74___block_34_tm_x;
_q___pip_5160_1_75___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___block_34_tm_x : _d___pip_5160_1_75___block_34_tm_x;
_q___pip_5160_1_76___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___block_34_tm_x : _d___pip_5160_1_76___block_34_tm_x;
_q___pip_5160_1_77___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___block_34_tm_x : _d___pip_5160_1_77___block_34_tm_x;
_q___pip_5160_1_78___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___block_34_tm_x : _d___pip_5160_1_78___block_34_tm_x;
_q___pip_5160_1_79___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___block_34_tm_x : _d___pip_5160_1_79___block_34_tm_x;
_q___pip_5160_1_80___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___block_34_tm_x : _d___pip_5160_1_80___block_34_tm_x;
_q___pip_5160_1_81___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___block_34_tm_x : _d___pip_5160_1_81___block_34_tm_x;
_q___pip_5160_1_82___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___block_34_tm_x : _d___pip_5160_1_82___block_34_tm_x;
_q___pip_5160_1_83___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___block_34_tm_x : _d___pip_5160_1_83___block_34_tm_x;
_q___pip_5160_1_84___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___block_34_tm_x : _d___pip_5160_1_84___block_34_tm_x;
_q___pip_5160_1_85___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___block_34_tm_x : _d___pip_5160_1_85___block_34_tm_x;
_q___pip_5160_1_86___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___block_34_tm_x : _d___pip_5160_1_86___block_34_tm_x;
_q___pip_5160_1_87___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___block_34_tm_x : _d___pip_5160_1_87___block_34_tm_x;
_q___pip_5160_1_88___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___block_34_tm_x : _d___pip_5160_1_88___block_34_tm_x;
_q___pip_5160_1_89___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___block_34_tm_x : _d___pip_5160_1_89___block_34_tm_x;
_q___pip_5160_1_90___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___block_34_tm_x : _d___pip_5160_1_90___block_34_tm_x;
_q___pip_5160_1_91___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___block_34_tm_x : _d___pip_5160_1_91___block_34_tm_x;
_q___pip_5160_1_92___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___block_34_tm_x : _d___pip_5160_1_92___block_34_tm_x;
_q___pip_5160_1_93___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___block_34_tm_x : _d___pip_5160_1_93___block_34_tm_x;
_q___pip_5160_1_94___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___block_34_tm_x : _d___pip_5160_1_94___block_34_tm_x;
_q___pip_5160_1_95___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___block_34_tm_x : _d___pip_5160_1_95___block_34_tm_x;
_q___pip_5160_1_96___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___block_34_tm_x : _d___pip_5160_1_96___block_34_tm_x;
_q___pip_5160_1_97___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___block_34_tm_x : _d___pip_5160_1_97___block_34_tm_x;
_q___pip_5160_1_98___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___block_34_tm_x : _d___pip_5160_1_98___block_34_tm_x;
_q___pip_5160_1_99___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___block_34_tm_x : _d___pip_5160_1_99___block_34_tm_x;
_q___pip_5160_1_100___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___block_34_tm_x : _d___pip_5160_1_100___block_34_tm_x;
_q___pip_5160_1_101___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___block_34_tm_x : _d___pip_5160_1_101___block_34_tm_x;
_q___pip_5160_1_102___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___block_34_tm_x : _d___pip_5160_1_102___block_34_tm_x;
_q___pip_5160_1_103___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___block_34_tm_x : _d___pip_5160_1_103___block_34_tm_x;
_q___pip_5160_1_104___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___block_34_tm_x : _d___pip_5160_1_104___block_34_tm_x;
_q___pip_5160_1_105___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___block_34_tm_x : _d___pip_5160_1_105___block_34_tm_x;
_q___pip_5160_1_106___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___block_34_tm_x : _d___pip_5160_1_106___block_34_tm_x;
_q___pip_5160_1_107___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___block_34_tm_x : _d___pip_5160_1_107___block_34_tm_x;
_q___pip_5160_1_108___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___block_34_tm_x : _d___pip_5160_1_108___block_34_tm_x;
_q___pip_5160_1_109___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___block_34_tm_x : _d___pip_5160_1_109___block_34_tm_x;
_q___pip_5160_1_110___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___block_34_tm_x : _d___pip_5160_1_110___block_34_tm_x;
_q___pip_5160_1_111___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___block_34_tm_x : _d___pip_5160_1_111___block_34_tm_x;
_q___pip_5160_1_112___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___block_34_tm_x : _d___pip_5160_1_112___block_34_tm_x;
_q___pip_5160_1_113___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___block_34_tm_x : _d___pip_5160_1_113___block_34_tm_x;
_q___pip_5160_1_114___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___block_34_tm_x : _d___pip_5160_1_114___block_34_tm_x;
_q___pip_5160_1_115___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___block_34_tm_x : _d___pip_5160_1_115___block_34_tm_x;
_q___pip_5160_1_116___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___block_34_tm_x : _d___pip_5160_1_116___block_34_tm_x;
_q___pip_5160_1_117___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___block_34_tm_x : _d___pip_5160_1_117___block_34_tm_x;
_q___pip_5160_1_118___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___block_34_tm_x : _d___pip_5160_1_118___block_34_tm_x;
_q___pip_5160_1_119___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___block_34_tm_x : _d___pip_5160_1_119___block_34_tm_x;
_q___pip_5160_1_120___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___block_34_tm_x : _d___pip_5160_1_120___block_34_tm_x;
_q___pip_5160_1_121___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___block_34_tm_x : _d___pip_5160_1_121___block_34_tm_x;
_q___pip_5160_1_122___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___block_34_tm_x : _d___pip_5160_1_122___block_34_tm_x;
_q___pip_5160_1_123___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___block_34_tm_x : _d___pip_5160_1_123___block_34_tm_x;
_q___pip_5160_1_124___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___block_34_tm_x : _d___pip_5160_1_124___block_34_tm_x;
_q___pip_5160_1_125___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___block_34_tm_x : _d___pip_5160_1_125___block_34_tm_x;
_q___pip_5160_1_126___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___block_34_tm_x : _d___pip_5160_1_126___block_34_tm_x;
_q___pip_5160_1_127___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___block_34_tm_x : _d___pip_5160_1_127___block_34_tm_x;
_q___pip_5160_1_128___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___block_34_tm_x : _d___pip_5160_1_128___block_34_tm_x;
_q___pip_5160_1_129___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___block_34_tm_x : _d___pip_5160_1_129___block_34_tm_x;
_q___pip_5160_1_130___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___block_34_tm_x : _d___pip_5160_1_130___block_34_tm_x;
_q___pip_5160_1_131___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___block_34_tm_x : _d___pip_5160_1_131___block_34_tm_x;
_q___pip_5160_1_132___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___block_34_tm_x : _d___pip_5160_1_132___block_34_tm_x;
_q___pip_5160_1_133___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___block_34_tm_x : _d___pip_5160_1_133___block_34_tm_x;
_q___pip_5160_1_134___block_34_tm_x <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___block_34_tm_x : _d___pip_5160_1_134___block_34_tm_x;
_q___pip_5160_1_6___block_34_tm_y <= _d___pip_5160_1_6___block_34_tm_y;
_q___pip_5160_1_7___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___block_34_tm_y : _d___pip_5160_1_7___block_34_tm_y;
_q___pip_5160_1_8___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___block_34_tm_y : _d___pip_5160_1_8___block_34_tm_y;
_q___pip_5160_1_9___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___block_34_tm_y : _d___pip_5160_1_9___block_34_tm_y;
_q___pip_5160_1_10___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___block_34_tm_y : _d___pip_5160_1_10___block_34_tm_y;
_q___pip_5160_1_11___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___block_34_tm_y : _d___pip_5160_1_11___block_34_tm_y;
_q___pip_5160_1_12___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___block_34_tm_y : _d___pip_5160_1_12___block_34_tm_y;
_q___pip_5160_1_13___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___block_34_tm_y : _d___pip_5160_1_13___block_34_tm_y;
_q___pip_5160_1_14___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___block_34_tm_y : _d___pip_5160_1_14___block_34_tm_y;
_q___pip_5160_1_15___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___block_34_tm_y : _d___pip_5160_1_15___block_34_tm_y;
_q___pip_5160_1_16___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___block_34_tm_y : _d___pip_5160_1_16___block_34_tm_y;
_q___pip_5160_1_17___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___block_34_tm_y : _d___pip_5160_1_17___block_34_tm_y;
_q___pip_5160_1_18___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___block_34_tm_y : _d___pip_5160_1_18___block_34_tm_y;
_q___pip_5160_1_19___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___block_34_tm_y : _d___pip_5160_1_19___block_34_tm_y;
_q___pip_5160_1_20___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___block_34_tm_y : _d___pip_5160_1_20___block_34_tm_y;
_q___pip_5160_1_21___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___block_34_tm_y : _d___pip_5160_1_21___block_34_tm_y;
_q___pip_5160_1_22___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___block_34_tm_y : _d___pip_5160_1_22___block_34_tm_y;
_q___pip_5160_1_23___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___block_34_tm_y : _d___pip_5160_1_23___block_34_tm_y;
_q___pip_5160_1_24___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___block_34_tm_y : _d___pip_5160_1_24___block_34_tm_y;
_q___pip_5160_1_25___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___block_34_tm_y : _d___pip_5160_1_25___block_34_tm_y;
_q___pip_5160_1_26___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___block_34_tm_y : _d___pip_5160_1_26___block_34_tm_y;
_q___pip_5160_1_27___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___block_34_tm_y : _d___pip_5160_1_27___block_34_tm_y;
_q___pip_5160_1_28___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___block_34_tm_y : _d___pip_5160_1_28___block_34_tm_y;
_q___pip_5160_1_29___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___block_34_tm_y : _d___pip_5160_1_29___block_34_tm_y;
_q___pip_5160_1_30___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___block_34_tm_y : _d___pip_5160_1_30___block_34_tm_y;
_q___pip_5160_1_31___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___block_34_tm_y : _d___pip_5160_1_31___block_34_tm_y;
_q___pip_5160_1_32___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___block_34_tm_y : _d___pip_5160_1_32___block_34_tm_y;
_q___pip_5160_1_33___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___block_34_tm_y : _d___pip_5160_1_33___block_34_tm_y;
_q___pip_5160_1_34___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___block_34_tm_y : _d___pip_5160_1_34___block_34_tm_y;
_q___pip_5160_1_35___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___block_34_tm_y : _d___pip_5160_1_35___block_34_tm_y;
_q___pip_5160_1_36___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___block_34_tm_y : _d___pip_5160_1_36___block_34_tm_y;
_q___pip_5160_1_37___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___block_34_tm_y : _d___pip_5160_1_37___block_34_tm_y;
_q___pip_5160_1_38___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___block_34_tm_y : _d___pip_5160_1_38___block_34_tm_y;
_q___pip_5160_1_39___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___block_34_tm_y : _d___pip_5160_1_39___block_34_tm_y;
_q___pip_5160_1_40___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___block_34_tm_y : _d___pip_5160_1_40___block_34_tm_y;
_q___pip_5160_1_41___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___block_34_tm_y : _d___pip_5160_1_41___block_34_tm_y;
_q___pip_5160_1_42___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___block_34_tm_y : _d___pip_5160_1_42___block_34_tm_y;
_q___pip_5160_1_43___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___block_34_tm_y : _d___pip_5160_1_43___block_34_tm_y;
_q___pip_5160_1_44___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___block_34_tm_y : _d___pip_5160_1_44___block_34_tm_y;
_q___pip_5160_1_45___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___block_34_tm_y : _d___pip_5160_1_45___block_34_tm_y;
_q___pip_5160_1_46___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___block_34_tm_y : _d___pip_5160_1_46___block_34_tm_y;
_q___pip_5160_1_47___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___block_34_tm_y : _d___pip_5160_1_47___block_34_tm_y;
_q___pip_5160_1_48___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___block_34_tm_y : _d___pip_5160_1_48___block_34_tm_y;
_q___pip_5160_1_49___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___block_34_tm_y : _d___pip_5160_1_49___block_34_tm_y;
_q___pip_5160_1_50___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___block_34_tm_y : _d___pip_5160_1_50___block_34_tm_y;
_q___pip_5160_1_51___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___block_34_tm_y : _d___pip_5160_1_51___block_34_tm_y;
_q___pip_5160_1_52___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___block_34_tm_y : _d___pip_5160_1_52___block_34_tm_y;
_q___pip_5160_1_53___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___block_34_tm_y : _d___pip_5160_1_53___block_34_tm_y;
_q___pip_5160_1_54___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___block_34_tm_y : _d___pip_5160_1_54___block_34_tm_y;
_q___pip_5160_1_55___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___block_34_tm_y : _d___pip_5160_1_55___block_34_tm_y;
_q___pip_5160_1_56___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___block_34_tm_y : _d___pip_5160_1_56___block_34_tm_y;
_q___pip_5160_1_57___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___block_34_tm_y : _d___pip_5160_1_57___block_34_tm_y;
_q___pip_5160_1_58___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___block_34_tm_y : _d___pip_5160_1_58___block_34_tm_y;
_q___pip_5160_1_59___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___block_34_tm_y : _d___pip_5160_1_59___block_34_tm_y;
_q___pip_5160_1_60___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___block_34_tm_y : _d___pip_5160_1_60___block_34_tm_y;
_q___pip_5160_1_61___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___block_34_tm_y : _d___pip_5160_1_61___block_34_tm_y;
_q___pip_5160_1_62___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___block_34_tm_y : _d___pip_5160_1_62___block_34_tm_y;
_q___pip_5160_1_63___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___block_34_tm_y : _d___pip_5160_1_63___block_34_tm_y;
_q___pip_5160_1_64___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___block_34_tm_y : _d___pip_5160_1_64___block_34_tm_y;
_q___pip_5160_1_65___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___block_34_tm_y : _d___pip_5160_1_65___block_34_tm_y;
_q___pip_5160_1_66___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___block_34_tm_y : _d___pip_5160_1_66___block_34_tm_y;
_q___pip_5160_1_67___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___block_34_tm_y : _d___pip_5160_1_67___block_34_tm_y;
_q___pip_5160_1_68___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___block_34_tm_y : _d___pip_5160_1_68___block_34_tm_y;
_q___pip_5160_1_69___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___block_34_tm_y : _d___pip_5160_1_69___block_34_tm_y;
_q___pip_5160_1_70___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___block_34_tm_y : _d___pip_5160_1_70___block_34_tm_y;
_q___pip_5160_1_71___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___block_34_tm_y : _d___pip_5160_1_71___block_34_tm_y;
_q___pip_5160_1_72___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___block_34_tm_y : _d___pip_5160_1_72___block_34_tm_y;
_q___pip_5160_1_73___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___block_34_tm_y : _d___pip_5160_1_73___block_34_tm_y;
_q___pip_5160_1_74___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___block_34_tm_y : _d___pip_5160_1_74___block_34_tm_y;
_q___pip_5160_1_75___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___block_34_tm_y : _d___pip_5160_1_75___block_34_tm_y;
_q___pip_5160_1_76___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___block_34_tm_y : _d___pip_5160_1_76___block_34_tm_y;
_q___pip_5160_1_77___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___block_34_tm_y : _d___pip_5160_1_77___block_34_tm_y;
_q___pip_5160_1_78___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___block_34_tm_y : _d___pip_5160_1_78___block_34_tm_y;
_q___pip_5160_1_79___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___block_34_tm_y : _d___pip_5160_1_79___block_34_tm_y;
_q___pip_5160_1_80___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___block_34_tm_y : _d___pip_5160_1_80___block_34_tm_y;
_q___pip_5160_1_81___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___block_34_tm_y : _d___pip_5160_1_81___block_34_tm_y;
_q___pip_5160_1_82___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___block_34_tm_y : _d___pip_5160_1_82___block_34_tm_y;
_q___pip_5160_1_83___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___block_34_tm_y : _d___pip_5160_1_83___block_34_tm_y;
_q___pip_5160_1_84___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___block_34_tm_y : _d___pip_5160_1_84___block_34_tm_y;
_q___pip_5160_1_85___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___block_34_tm_y : _d___pip_5160_1_85___block_34_tm_y;
_q___pip_5160_1_86___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___block_34_tm_y : _d___pip_5160_1_86___block_34_tm_y;
_q___pip_5160_1_87___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___block_34_tm_y : _d___pip_5160_1_87___block_34_tm_y;
_q___pip_5160_1_88___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___block_34_tm_y : _d___pip_5160_1_88___block_34_tm_y;
_q___pip_5160_1_89___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___block_34_tm_y : _d___pip_5160_1_89___block_34_tm_y;
_q___pip_5160_1_90___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___block_34_tm_y : _d___pip_5160_1_90___block_34_tm_y;
_q___pip_5160_1_91___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___block_34_tm_y : _d___pip_5160_1_91___block_34_tm_y;
_q___pip_5160_1_92___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___block_34_tm_y : _d___pip_5160_1_92___block_34_tm_y;
_q___pip_5160_1_93___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___block_34_tm_y : _d___pip_5160_1_93___block_34_tm_y;
_q___pip_5160_1_94___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___block_34_tm_y : _d___pip_5160_1_94___block_34_tm_y;
_q___pip_5160_1_95___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___block_34_tm_y : _d___pip_5160_1_95___block_34_tm_y;
_q___pip_5160_1_96___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___block_34_tm_y : _d___pip_5160_1_96___block_34_tm_y;
_q___pip_5160_1_97___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___block_34_tm_y : _d___pip_5160_1_97___block_34_tm_y;
_q___pip_5160_1_98___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___block_34_tm_y : _d___pip_5160_1_98___block_34_tm_y;
_q___pip_5160_1_99___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___block_34_tm_y : _d___pip_5160_1_99___block_34_tm_y;
_q___pip_5160_1_100___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___block_34_tm_y : _d___pip_5160_1_100___block_34_tm_y;
_q___pip_5160_1_101___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___block_34_tm_y : _d___pip_5160_1_101___block_34_tm_y;
_q___pip_5160_1_102___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___block_34_tm_y : _d___pip_5160_1_102___block_34_tm_y;
_q___pip_5160_1_103___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___block_34_tm_y : _d___pip_5160_1_103___block_34_tm_y;
_q___pip_5160_1_104___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___block_34_tm_y : _d___pip_5160_1_104___block_34_tm_y;
_q___pip_5160_1_105___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___block_34_tm_y : _d___pip_5160_1_105___block_34_tm_y;
_q___pip_5160_1_106___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___block_34_tm_y : _d___pip_5160_1_106___block_34_tm_y;
_q___pip_5160_1_107___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___block_34_tm_y : _d___pip_5160_1_107___block_34_tm_y;
_q___pip_5160_1_108___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___block_34_tm_y : _d___pip_5160_1_108___block_34_tm_y;
_q___pip_5160_1_109___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___block_34_tm_y : _d___pip_5160_1_109___block_34_tm_y;
_q___pip_5160_1_110___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___block_34_tm_y : _d___pip_5160_1_110___block_34_tm_y;
_q___pip_5160_1_111___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___block_34_tm_y : _d___pip_5160_1_111___block_34_tm_y;
_q___pip_5160_1_112___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___block_34_tm_y : _d___pip_5160_1_112___block_34_tm_y;
_q___pip_5160_1_113___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___block_34_tm_y : _d___pip_5160_1_113___block_34_tm_y;
_q___pip_5160_1_114___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___block_34_tm_y : _d___pip_5160_1_114___block_34_tm_y;
_q___pip_5160_1_115___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___block_34_tm_y : _d___pip_5160_1_115___block_34_tm_y;
_q___pip_5160_1_116___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___block_34_tm_y : _d___pip_5160_1_116___block_34_tm_y;
_q___pip_5160_1_117___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___block_34_tm_y : _d___pip_5160_1_117___block_34_tm_y;
_q___pip_5160_1_118___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___block_34_tm_y : _d___pip_5160_1_118___block_34_tm_y;
_q___pip_5160_1_119___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___block_34_tm_y : _d___pip_5160_1_119___block_34_tm_y;
_q___pip_5160_1_120___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___block_34_tm_y : _d___pip_5160_1_120___block_34_tm_y;
_q___pip_5160_1_121___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___block_34_tm_y : _d___pip_5160_1_121___block_34_tm_y;
_q___pip_5160_1_122___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___block_34_tm_y : _d___pip_5160_1_122___block_34_tm_y;
_q___pip_5160_1_123___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___block_34_tm_y : _d___pip_5160_1_123___block_34_tm_y;
_q___pip_5160_1_124___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___block_34_tm_y : _d___pip_5160_1_124___block_34_tm_y;
_q___pip_5160_1_125___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___block_34_tm_y : _d___pip_5160_1_125___block_34_tm_y;
_q___pip_5160_1_126___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___block_34_tm_y : _d___pip_5160_1_126___block_34_tm_y;
_q___pip_5160_1_127___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___block_34_tm_y : _d___pip_5160_1_127___block_34_tm_y;
_q___pip_5160_1_128___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___block_34_tm_y : _d___pip_5160_1_128___block_34_tm_y;
_q___pip_5160_1_129___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___block_34_tm_y : _d___pip_5160_1_129___block_34_tm_y;
_q___pip_5160_1_130___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___block_34_tm_y : _d___pip_5160_1_130___block_34_tm_y;
_q___pip_5160_1_131___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___block_34_tm_y : _d___pip_5160_1_131___block_34_tm_y;
_q___pip_5160_1_132___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___block_34_tm_y : _d___pip_5160_1_132___block_34_tm_y;
_q___pip_5160_1_133___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___block_34_tm_y : _d___pip_5160_1_133___block_34_tm_y;
_q___pip_5160_1_134___block_34_tm_y <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___block_34_tm_y : _d___pip_5160_1_134___block_34_tm_y;
_q___pip_5160_1_6___block_34_tm_z <= _d___pip_5160_1_6___block_34_tm_z;
_q___pip_5160_1_7___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___block_34_tm_z : _d___pip_5160_1_7___block_34_tm_z;
_q___pip_5160_1_8___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___block_34_tm_z : _d___pip_5160_1_8___block_34_tm_z;
_q___pip_5160_1_9___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___block_34_tm_z : _d___pip_5160_1_9___block_34_tm_z;
_q___pip_5160_1_10___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___block_34_tm_z : _d___pip_5160_1_10___block_34_tm_z;
_q___pip_5160_1_11___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___block_34_tm_z : _d___pip_5160_1_11___block_34_tm_z;
_q___pip_5160_1_12___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___block_34_tm_z : _d___pip_5160_1_12___block_34_tm_z;
_q___pip_5160_1_13___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___block_34_tm_z : _d___pip_5160_1_13___block_34_tm_z;
_q___pip_5160_1_14___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___block_34_tm_z : _d___pip_5160_1_14___block_34_tm_z;
_q___pip_5160_1_15___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___block_34_tm_z : _d___pip_5160_1_15___block_34_tm_z;
_q___pip_5160_1_16___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___block_34_tm_z : _d___pip_5160_1_16___block_34_tm_z;
_q___pip_5160_1_17___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___block_34_tm_z : _d___pip_5160_1_17___block_34_tm_z;
_q___pip_5160_1_18___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___block_34_tm_z : _d___pip_5160_1_18___block_34_tm_z;
_q___pip_5160_1_19___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___block_34_tm_z : _d___pip_5160_1_19___block_34_tm_z;
_q___pip_5160_1_20___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___block_34_tm_z : _d___pip_5160_1_20___block_34_tm_z;
_q___pip_5160_1_21___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___block_34_tm_z : _d___pip_5160_1_21___block_34_tm_z;
_q___pip_5160_1_22___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___block_34_tm_z : _d___pip_5160_1_22___block_34_tm_z;
_q___pip_5160_1_23___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___block_34_tm_z : _d___pip_5160_1_23___block_34_tm_z;
_q___pip_5160_1_24___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___block_34_tm_z : _d___pip_5160_1_24___block_34_tm_z;
_q___pip_5160_1_25___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___block_34_tm_z : _d___pip_5160_1_25___block_34_tm_z;
_q___pip_5160_1_26___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___block_34_tm_z : _d___pip_5160_1_26___block_34_tm_z;
_q___pip_5160_1_27___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___block_34_tm_z : _d___pip_5160_1_27___block_34_tm_z;
_q___pip_5160_1_28___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___block_34_tm_z : _d___pip_5160_1_28___block_34_tm_z;
_q___pip_5160_1_29___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___block_34_tm_z : _d___pip_5160_1_29___block_34_tm_z;
_q___pip_5160_1_30___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___block_34_tm_z : _d___pip_5160_1_30___block_34_tm_z;
_q___pip_5160_1_31___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___block_34_tm_z : _d___pip_5160_1_31___block_34_tm_z;
_q___pip_5160_1_32___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___block_34_tm_z : _d___pip_5160_1_32___block_34_tm_z;
_q___pip_5160_1_33___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___block_34_tm_z : _d___pip_5160_1_33___block_34_tm_z;
_q___pip_5160_1_34___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___block_34_tm_z : _d___pip_5160_1_34___block_34_tm_z;
_q___pip_5160_1_35___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___block_34_tm_z : _d___pip_5160_1_35___block_34_tm_z;
_q___pip_5160_1_36___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___block_34_tm_z : _d___pip_5160_1_36___block_34_tm_z;
_q___pip_5160_1_37___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___block_34_tm_z : _d___pip_5160_1_37___block_34_tm_z;
_q___pip_5160_1_38___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___block_34_tm_z : _d___pip_5160_1_38___block_34_tm_z;
_q___pip_5160_1_39___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___block_34_tm_z : _d___pip_5160_1_39___block_34_tm_z;
_q___pip_5160_1_40___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___block_34_tm_z : _d___pip_5160_1_40___block_34_tm_z;
_q___pip_5160_1_41___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___block_34_tm_z : _d___pip_5160_1_41___block_34_tm_z;
_q___pip_5160_1_42___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___block_34_tm_z : _d___pip_5160_1_42___block_34_tm_z;
_q___pip_5160_1_43___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___block_34_tm_z : _d___pip_5160_1_43___block_34_tm_z;
_q___pip_5160_1_44___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___block_34_tm_z : _d___pip_5160_1_44___block_34_tm_z;
_q___pip_5160_1_45___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___block_34_tm_z : _d___pip_5160_1_45___block_34_tm_z;
_q___pip_5160_1_46___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___block_34_tm_z : _d___pip_5160_1_46___block_34_tm_z;
_q___pip_5160_1_47___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___block_34_tm_z : _d___pip_5160_1_47___block_34_tm_z;
_q___pip_5160_1_48___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___block_34_tm_z : _d___pip_5160_1_48___block_34_tm_z;
_q___pip_5160_1_49___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___block_34_tm_z : _d___pip_5160_1_49___block_34_tm_z;
_q___pip_5160_1_50___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___block_34_tm_z : _d___pip_5160_1_50___block_34_tm_z;
_q___pip_5160_1_51___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___block_34_tm_z : _d___pip_5160_1_51___block_34_tm_z;
_q___pip_5160_1_52___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___block_34_tm_z : _d___pip_5160_1_52___block_34_tm_z;
_q___pip_5160_1_53___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___block_34_tm_z : _d___pip_5160_1_53___block_34_tm_z;
_q___pip_5160_1_54___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___block_34_tm_z : _d___pip_5160_1_54___block_34_tm_z;
_q___pip_5160_1_55___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___block_34_tm_z : _d___pip_5160_1_55___block_34_tm_z;
_q___pip_5160_1_56___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___block_34_tm_z : _d___pip_5160_1_56___block_34_tm_z;
_q___pip_5160_1_57___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___block_34_tm_z : _d___pip_5160_1_57___block_34_tm_z;
_q___pip_5160_1_58___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___block_34_tm_z : _d___pip_5160_1_58___block_34_tm_z;
_q___pip_5160_1_59___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___block_34_tm_z : _d___pip_5160_1_59___block_34_tm_z;
_q___pip_5160_1_60___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___block_34_tm_z : _d___pip_5160_1_60___block_34_tm_z;
_q___pip_5160_1_61___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___block_34_tm_z : _d___pip_5160_1_61___block_34_tm_z;
_q___pip_5160_1_62___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___block_34_tm_z : _d___pip_5160_1_62___block_34_tm_z;
_q___pip_5160_1_63___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___block_34_tm_z : _d___pip_5160_1_63___block_34_tm_z;
_q___pip_5160_1_64___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___block_34_tm_z : _d___pip_5160_1_64___block_34_tm_z;
_q___pip_5160_1_65___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___block_34_tm_z : _d___pip_5160_1_65___block_34_tm_z;
_q___pip_5160_1_66___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___block_34_tm_z : _d___pip_5160_1_66___block_34_tm_z;
_q___pip_5160_1_67___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___block_34_tm_z : _d___pip_5160_1_67___block_34_tm_z;
_q___pip_5160_1_68___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___block_34_tm_z : _d___pip_5160_1_68___block_34_tm_z;
_q___pip_5160_1_69___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___block_34_tm_z : _d___pip_5160_1_69___block_34_tm_z;
_q___pip_5160_1_70___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___block_34_tm_z : _d___pip_5160_1_70___block_34_tm_z;
_q___pip_5160_1_71___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___block_34_tm_z : _d___pip_5160_1_71___block_34_tm_z;
_q___pip_5160_1_72___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___block_34_tm_z : _d___pip_5160_1_72___block_34_tm_z;
_q___pip_5160_1_73___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___block_34_tm_z : _d___pip_5160_1_73___block_34_tm_z;
_q___pip_5160_1_74___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___block_34_tm_z : _d___pip_5160_1_74___block_34_tm_z;
_q___pip_5160_1_75___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___block_34_tm_z : _d___pip_5160_1_75___block_34_tm_z;
_q___pip_5160_1_76___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___block_34_tm_z : _d___pip_5160_1_76___block_34_tm_z;
_q___pip_5160_1_77___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___block_34_tm_z : _d___pip_5160_1_77___block_34_tm_z;
_q___pip_5160_1_78___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___block_34_tm_z : _d___pip_5160_1_78___block_34_tm_z;
_q___pip_5160_1_79___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___block_34_tm_z : _d___pip_5160_1_79___block_34_tm_z;
_q___pip_5160_1_80___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___block_34_tm_z : _d___pip_5160_1_80___block_34_tm_z;
_q___pip_5160_1_81___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___block_34_tm_z : _d___pip_5160_1_81___block_34_tm_z;
_q___pip_5160_1_82___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___block_34_tm_z : _d___pip_5160_1_82___block_34_tm_z;
_q___pip_5160_1_83___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___block_34_tm_z : _d___pip_5160_1_83___block_34_tm_z;
_q___pip_5160_1_84___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___block_34_tm_z : _d___pip_5160_1_84___block_34_tm_z;
_q___pip_5160_1_85___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___block_34_tm_z : _d___pip_5160_1_85___block_34_tm_z;
_q___pip_5160_1_86___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___block_34_tm_z : _d___pip_5160_1_86___block_34_tm_z;
_q___pip_5160_1_87___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___block_34_tm_z : _d___pip_5160_1_87___block_34_tm_z;
_q___pip_5160_1_88___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___block_34_tm_z : _d___pip_5160_1_88___block_34_tm_z;
_q___pip_5160_1_89___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___block_34_tm_z : _d___pip_5160_1_89___block_34_tm_z;
_q___pip_5160_1_90___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___block_34_tm_z : _d___pip_5160_1_90___block_34_tm_z;
_q___pip_5160_1_91___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___block_34_tm_z : _d___pip_5160_1_91___block_34_tm_z;
_q___pip_5160_1_92___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___block_34_tm_z : _d___pip_5160_1_92___block_34_tm_z;
_q___pip_5160_1_93___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___block_34_tm_z : _d___pip_5160_1_93___block_34_tm_z;
_q___pip_5160_1_94___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___block_34_tm_z : _d___pip_5160_1_94___block_34_tm_z;
_q___pip_5160_1_95___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___block_34_tm_z : _d___pip_5160_1_95___block_34_tm_z;
_q___pip_5160_1_96___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___block_34_tm_z : _d___pip_5160_1_96___block_34_tm_z;
_q___pip_5160_1_97___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___block_34_tm_z : _d___pip_5160_1_97___block_34_tm_z;
_q___pip_5160_1_98___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___block_34_tm_z : _d___pip_5160_1_98___block_34_tm_z;
_q___pip_5160_1_99___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___block_34_tm_z : _d___pip_5160_1_99___block_34_tm_z;
_q___pip_5160_1_100___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___block_34_tm_z : _d___pip_5160_1_100___block_34_tm_z;
_q___pip_5160_1_101___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___block_34_tm_z : _d___pip_5160_1_101___block_34_tm_z;
_q___pip_5160_1_102___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___block_34_tm_z : _d___pip_5160_1_102___block_34_tm_z;
_q___pip_5160_1_103___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___block_34_tm_z : _d___pip_5160_1_103___block_34_tm_z;
_q___pip_5160_1_104___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___block_34_tm_z : _d___pip_5160_1_104___block_34_tm_z;
_q___pip_5160_1_105___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___block_34_tm_z : _d___pip_5160_1_105___block_34_tm_z;
_q___pip_5160_1_106___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___block_34_tm_z : _d___pip_5160_1_106___block_34_tm_z;
_q___pip_5160_1_107___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___block_34_tm_z : _d___pip_5160_1_107___block_34_tm_z;
_q___pip_5160_1_108___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___block_34_tm_z : _d___pip_5160_1_108___block_34_tm_z;
_q___pip_5160_1_109___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___block_34_tm_z : _d___pip_5160_1_109___block_34_tm_z;
_q___pip_5160_1_110___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___block_34_tm_z : _d___pip_5160_1_110___block_34_tm_z;
_q___pip_5160_1_111___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___block_34_tm_z : _d___pip_5160_1_111___block_34_tm_z;
_q___pip_5160_1_112___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___block_34_tm_z : _d___pip_5160_1_112___block_34_tm_z;
_q___pip_5160_1_113___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___block_34_tm_z : _d___pip_5160_1_113___block_34_tm_z;
_q___pip_5160_1_114___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___block_34_tm_z : _d___pip_5160_1_114___block_34_tm_z;
_q___pip_5160_1_115___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___block_34_tm_z : _d___pip_5160_1_115___block_34_tm_z;
_q___pip_5160_1_116___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___block_34_tm_z : _d___pip_5160_1_116___block_34_tm_z;
_q___pip_5160_1_117___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___block_34_tm_z : _d___pip_5160_1_117___block_34_tm_z;
_q___pip_5160_1_118___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___block_34_tm_z : _d___pip_5160_1_118___block_34_tm_z;
_q___pip_5160_1_119___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___block_34_tm_z : _d___pip_5160_1_119___block_34_tm_z;
_q___pip_5160_1_120___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___block_34_tm_z : _d___pip_5160_1_120___block_34_tm_z;
_q___pip_5160_1_121___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___block_34_tm_z : _d___pip_5160_1_121___block_34_tm_z;
_q___pip_5160_1_122___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___block_34_tm_z : _d___pip_5160_1_122___block_34_tm_z;
_q___pip_5160_1_123___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___block_34_tm_z : _d___pip_5160_1_123___block_34_tm_z;
_q___pip_5160_1_124___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___block_34_tm_z : _d___pip_5160_1_124___block_34_tm_z;
_q___pip_5160_1_125___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___block_34_tm_z : _d___pip_5160_1_125___block_34_tm_z;
_q___pip_5160_1_126___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___block_34_tm_z : _d___pip_5160_1_126___block_34_tm_z;
_q___pip_5160_1_127___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___block_34_tm_z : _d___pip_5160_1_127___block_34_tm_z;
_q___pip_5160_1_128___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___block_34_tm_z : _d___pip_5160_1_128___block_34_tm_z;
_q___pip_5160_1_129___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___block_34_tm_z : _d___pip_5160_1_129___block_34_tm_z;
_q___pip_5160_1_130___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___block_34_tm_z : _d___pip_5160_1_130___block_34_tm_z;
_q___pip_5160_1_131___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___block_34_tm_z : _d___pip_5160_1_131___block_34_tm_z;
_q___pip_5160_1_132___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___block_34_tm_z : _d___pip_5160_1_132___block_34_tm_z;
_q___pip_5160_1_133___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___block_34_tm_z : _d___pip_5160_1_133___block_34_tm_z;
_q___pip_5160_1_134___block_34_tm_z <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___block_34_tm_z : _d___pip_5160_1_134___block_34_tm_z;
_q___pip_5160_1_6___block_40_dt_x <= _d___pip_5160_1_6___block_40_dt_x;
_q___pip_5160_1_7___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___block_40_dt_x : _d___pip_5160_1_7___block_40_dt_x;
_q___pip_5160_1_8___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___block_40_dt_x : _d___pip_5160_1_8___block_40_dt_x;
_q___pip_5160_1_9___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___block_40_dt_x : _d___pip_5160_1_9___block_40_dt_x;
_q___pip_5160_1_10___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___block_40_dt_x : _d___pip_5160_1_10___block_40_dt_x;
_q___pip_5160_1_11___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___block_40_dt_x : _d___pip_5160_1_11___block_40_dt_x;
_q___pip_5160_1_12___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___block_40_dt_x : _d___pip_5160_1_12___block_40_dt_x;
_q___pip_5160_1_13___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___block_40_dt_x : _d___pip_5160_1_13___block_40_dt_x;
_q___pip_5160_1_14___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___block_40_dt_x : _d___pip_5160_1_14___block_40_dt_x;
_q___pip_5160_1_15___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___block_40_dt_x : _d___pip_5160_1_15___block_40_dt_x;
_q___pip_5160_1_16___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___block_40_dt_x : _d___pip_5160_1_16___block_40_dt_x;
_q___pip_5160_1_17___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___block_40_dt_x : _d___pip_5160_1_17___block_40_dt_x;
_q___pip_5160_1_18___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___block_40_dt_x : _d___pip_5160_1_18___block_40_dt_x;
_q___pip_5160_1_19___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___block_40_dt_x : _d___pip_5160_1_19___block_40_dt_x;
_q___pip_5160_1_20___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___block_40_dt_x : _d___pip_5160_1_20___block_40_dt_x;
_q___pip_5160_1_21___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___block_40_dt_x : _d___pip_5160_1_21___block_40_dt_x;
_q___pip_5160_1_22___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___block_40_dt_x : _d___pip_5160_1_22___block_40_dt_x;
_q___pip_5160_1_23___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___block_40_dt_x : _d___pip_5160_1_23___block_40_dt_x;
_q___pip_5160_1_24___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___block_40_dt_x : _d___pip_5160_1_24___block_40_dt_x;
_q___pip_5160_1_25___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___block_40_dt_x : _d___pip_5160_1_25___block_40_dt_x;
_q___pip_5160_1_26___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___block_40_dt_x : _d___pip_5160_1_26___block_40_dt_x;
_q___pip_5160_1_27___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___block_40_dt_x : _d___pip_5160_1_27___block_40_dt_x;
_q___pip_5160_1_28___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___block_40_dt_x : _d___pip_5160_1_28___block_40_dt_x;
_q___pip_5160_1_29___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___block_40_dt_x : _d___pip_5160_1_29___block_40_dt_x;
_q___pip_5160_1_30___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___block_40_dt_x : _d___pip_5160_1_30___block_40_dt_x;
_q___pip_5160_1_31___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___block_40_dt_x : _d___pip_5160_1_31___block_40_dt_x;
_q___pip_5160_1_32___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___block_40_dt_x : _d___pip_5160_1_32___block_40_dt_x;
_q___pip_5160_1_33___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___block_40_dt_x : _d___pip_5160_1_33___block_40_dt_x;
_q___pip_5160_1_34___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___block_40_dt_x : _d___pip_5160_1_34___block_40_dt_x;
_q___pip_5160_1_35___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___block_40_dt_x : _d___pip_5160_1_35___block_40_dt_x;
_q___pip_5160_1_36___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___block_40_dt_x : _d___pip_5160_1_36___block_40_dt_x;
_q___pip_5160_1_37___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___block_40_dt_x : _d___pip_5160_1_37___block_40_dt_x;
_q___pip_5160_1_38___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___block_40_dt_x : _d___pip_5160_1_38___block_40_dt_x;
_q___pip_5160_1_39___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___block_40_dt_x : _d___pip_5160_1_39___block_40_dt_x;
_q___pip_5160_1_40___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___block_40_dt_x : _d___pip_5160_1_40___block_40_dt_x;
_q___pip_5160_1_41___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___block_40_dt_x : _d___pip_5160_1_41___block_40_dt_x;
_q___pip_5160_1_42___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___block_40_dt_x : _d___pip_5160_1_42___block_40_dt_x;
_q___pip_5160_1_43___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___block_40_dt_x : _d___pip_5160_1_43___block_40_dt_x;
_q___pip_5160_1_44___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___block_40_dt_x : _d___pip_5160_1_44___block_40_dt_x;
_q___pip_5160_1_45___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___block_40_dt_x : _d___pip_5160_1_45___block_40_dt_x;
_q___pip_5160_1_46___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___block_40_dt_x : _d___pip_5160_1_46___block_40_dt_x;
_q___pip_5160_1_47___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___block_40_dt_x : _d___pip_5160_1_47___block_40_dt_x;
_q___pip_5160_1_48___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___block_40_dt_x : _d___pip_5160_1_48___block_40_dt_x;
_q___pip_5160_1_49___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___block_40_dt_x : _d___pip_5160_1_49___block_40_dt_x;
_q___pip_5160_1_50___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___block_40_dt_x : _d___pip_5160_1_50___block_40_dt_x;
_q___pip_5160_1_51___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___block_40_dt_x : _d___pip_5160_1_51___block_40_dt_x;
_q___pip_5160_1_52___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___block_40_dt_x : _d___pip_5160_1_52___block_40_dt_x;
_q___pip_5160_1_53___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___block_40_dt_x : _d___pip_5160_1_53___block_40_dt_x;
_q___pip_5160_1_54___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___block_40_dt_x : _d___pip_5160_1_54___block_40_dt_x;
_q___pip_5160_1_55___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___block_40_dt_x : _d___pip_5160_1_55___block_40_dt_x;
_q___pip_5160_1_56___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___block_40_dt_x : _d___pip_5160_1_56___block_40_dt_x;
_q___pip_5160_1_57___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___block_40_dt_x : _d___pip_5160_1_57___block_40_dt_x;
_q___pip_5160_1_58___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___block_40_dt_x : _d___pip_5160_1_58___block_40_dt_x;
_q___pip_5160_1_59___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___block_40_dt_x : _d___pip_5160_1_59___block_40_dt_x;
_q___pip_5160_1_60___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___block_40_dt_x : _d___pip_5160_1_60___block_40_dt_x;
_q___pip_5160_1_61___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___block_40_dt_x : _d___pip_5160_1_61___block_40_dt_x;
_q___pip_5160_1_62___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___block_40_dt_x : _d___pip_5160_1_62___block_40_dt_x;
_q___pip_5160_1_63___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___block_40_dt_x : _d___pip_5160_1_63___block_40_dt_x;
_q___pip_5160_1_64___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___block_40_dt_x : _d___pip_5160_1_64___block_40_dt_x;
_q___pip_5160_1_65___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___block_40_dt_x : _d___pip_5160_1_65___block_40_dt_x;
_q___pip_5160_1_66___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___block_40_dt_x : _d___pip_5160_1_66___block_40_dt_x;
_q___pip_5160_1_67___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___block_40_dt_x : _d___pip_5160_1_67___block_40_dt_x;
_q___pip_5160_1_68___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___block_40_dt_x : _d___pip_5160_1_68___block_40_dt_x;
_q___pip_5160_1_69___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___block_40_dt_x : _d___pip_5160_1_69___block_40_dt_x;
_q___pip_5160_1_70___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___block_40_dt_x : _d___pip_5160_1_70___block_40_dt_x;
_q___pip_5160_1_71___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___block_40_dt_x : _d___pip_5160_1_71___block_40_dt_x;
_q___pip_5160_1_72___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___block_40_dt_x : _d___pip_5160_1_72___block_40_dt_x;
_q___pip_5160_1_73___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___block_40_dt_x : _d___pip_5160_1_73___block_40_dt_x;
_q___pip_5160_1_74___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___block_40_dt_x : _d___pip_5160_1_74___block_40_dt_x;
_q___pip_5160_1_75___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___block_40_dt_x : _d___pip_5160_1_75___block_40_dt_x;
_q___pip_5160_1_76___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___block_40_dt_x : _d___pip_5160_1_76___block_40_dt_x;
_q___pip_5160_1_77___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___block_40_dt_x : _d___pip_5160_1_77___block_40_dt_x;
_q___pip_5160_1_78___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___block_40_dt_x : _d___pip_5160_1_78___block_40_dt_x;
_q___pip_5160_1_79___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___block_40_dt_x : _d___pip_5160_1_79___block_40_dt_x;
_q___pip_5160_1_80___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___block_40_dt_x : _d___pip_5160_1_80___block_40_dt_x;
_q___pip_5160_1_81___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___block_40_dt_x : _d___pip_5160_1_81___block_40_dt_x;
_q___pip_5160_1_82___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___block_40_dt_x : _d___pip_5160_1_82___block_40_dt_x;
_q___pip_5160_1_83___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___block_40_dt_x : _d___pip_5160_1_83___block_40_dt_x;
_q___pip_5160_1_84___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___block_40_dt_x : _d___pip_5160_1_84___block_40_dt_x;
_q___pip_5160_1_85___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___block_40_dt_x : _d___pip_5160_1_85___block_40_dt_x;
_q___pip_5160_1_86___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___block_40_dt_x : _d___pip_5160_1_86___block_40_dt_x;
_q___pip_5160_1_87___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___block_40_dt_x : _d___pip_5160_1_87___block_40_dt_x;
_q___pip_5160_1_88___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___block_40_dt_x : _d___pip_5160_1_88___block_40_dt_x;
_q___pip_5160_1_89___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___block_40_dt_x : _d___pip_5160_1_89___block_40_dt_x;
_q___pip_5160_1_90___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___block_40_dt_x : _d___pip_5160_1_90___block_40_dt_x;
_q___pip_5160_1_91___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___block_40_dt_x : _d___pip_5160_1_91___block_40_dt_x;
_q___pip_5160_1_92___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___block_40_dt_x : _d___pip_5160_1_92___block_40_dt_x;
_q___pip_5160_1_93___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___block_40_dt_x : _d___pip_5160_1_93___block_40_dt_x;
_q___pip_5160_1_94___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___block_40_dt_x : _d___pip_5160_1_94___block_40_dt_x;
_q___pip_5160_1_95___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___block_40_dt_x : _d___pip_5160_1_95___block_40_dt_x;
_q___pip_5160_1_96___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___block_40_dt_x : _d___pip_5160_1_96___block_40_dt_x;
_q___pip_5160_1_97___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___block_40_dt_x : _d___pip_5160_1_97___block_40_dt_x;
_q___pip_5160_1_98___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___block_40_dt_x : _d___pip_5160_1_98___block_40_dt_x;
_q___pip_5160_1_99___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___block_40_dt_x : _d___pip_5160_1_99___block_40_dt_x;
_q___pip_5160_1_100___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___block_40_dt_x : _d___pip_5160_1_100___block_40_dt_x;
_q___pip_5160_1_101___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___block_40_dt_x : _d___pip_5160_1_101___block_40_dt_x;
_q___pip_5160_1_102___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___block_40_dt_x : _d___pip_5160_1_102___block_40_dt_x;
_q___pip_5160_1_103___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___block_40_dt_x : _d___pip_5160_1_103___block_40_dt_x;
_q___pip_5160_1_104___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___block_40_dt_x : _d___pip_5160_1_104___block_40_dt_x;
_q___pip_5160_1_105___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___block_40_dt_x : _d___pip_5160_1_105___block_40_dt_x;
_q___pip_5160_1_106___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___block_40_dt_x : _d___pip_5160_1_106___block_40_dt_x;
_q___pip_5160_1_107___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___block_40_dt_x : _d___pip_5160_1_107___block_40_dt_x;
_q___pip_5160_1_108___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___block_40_dt_x : _d___pip_5160_1_108___block_40_dt_x;
_q___pip_5160_1_109___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___block_40_dt_x : _d___pip_5160_1_109___block_40_dt_x;
_q___pip_5160_1_110___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___block_40_dt_x : _d___pip_5160_1_110___block_40_dt_x;
_q___pip_5160_1_111___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___block_40_dt_x : _d___pip_5160_1_111___block_40_dt_x;
_q___pip_5160_1_112___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___block_40_dt_x : _d___pip_5160_1_112___block_40_dt_x;
_q___pip_5160_1_113___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___block_40_dt_x : _d___pip_5160_1_113___block_40_dt_x;
_q___pip_5160_1_114___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___block_40_dt_x : _d___pip_5160_1_114___block_40_dt_x;
_q___pip_5160_1_115___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___block_40_dt_x : _d___pip_5160_1_115___block_40_dt_x;
_q___pip_5160_1_116___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___block_40_dt_x : _d___pip_5160_1_116___block_40_dt_x;
_q___pip_5160_1_117___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___block_40_dt_x : _d___pip_5160_1_117___block_40_dt_x;
_q___pip_5160_1_118___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___block_40_dt_x : _d___pip_5160_1_118___block_40_dt_x;
_q___pip_5160_1_119___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___block_40_dt_x : _d___pip_5160_1_119___block_40_dt_x;
_q___pip_5160_1_120___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___block_40_dt_x : _d___pip_5160_1_120___block_40_dt_x;
_q___pip_5160_1_121___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___block_40_dt_x : _d___pip_5160_1_121___block_40_dt_x;
_q___pip_5160_1_122___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___block_40_dt_x : _d___pip_5160_1_122___block_40_dt_x;
_q___pip_5160_1_123___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___block_40_dt_x : _d___pip_5160_1_123___block_40_dt_x;
_q___pip_5160_1_124___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___block_40_dt_x : _d___pip_5160_1_124___block_40_dt_x;
_q___pip_5160_1_125___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___block_40_dt_x : _d___pip_5160_1_125___block_40_dt_x;
_q___pip_5160_1_126___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___block_40_dt_x : _d___pip_5160_1_126___block_40_dt_x;
_q___pip_5160_1_127___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___block_40_dt_x : _d___pip_5160_1_127___block_40_dt_x;
_q___pip_5160_1_128___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___block_40_dt_x : _d___pip_5160_1_128___block_40_dt_x;
_q___pip_5160_1_129___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___block_40_dt_x : _d___pip_5160_1_129___block_40_dt_x;
_q___pip_5160_1_130___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___block_40_dt_x : _d___pip_5160_1_130___block_40_dt_x;
_q___pip_5160_1_131___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___block_40_dt_x : _d___pip_5160_1_131___block_40_dt_x;
_q___pip_5160_1_132___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___block_40_dt_x : _d___pip_5160_1_132___block_40_dt_x;
_q___pip_5160_1_133___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___block_40_dt_x : _d___pip_5160_1_133___block_40_dt_x;
_q___pip_5160_1_134___block_40_dt_x <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___block_40_dt_x : _d___pip_5160_1_134___block_40_dt_x;
_q___pip_5160_1_6___block_40_dt_y <= _d___pip_5160_1_6___block_40_dt_y;
_q___pip_5160_1_7___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___block_40_dt_y : _d___pip_5160_1_7___block_40_dt_y;
_q___pip_5160_1_8___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___block_40_dt_y : _d___pip_5160_1_8___block_40_dt_y;
_q___pip_5160_1_9___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___block_40_dt_y : _d___pip_5160_1_9___block_40_dt_y;
_q___pip_5160_1_10___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___block_40_dt_y : _d___pip_5160_1_10___block_40_dt_y;
_q___pip_5160_1_11___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___block_40_dt_y : _d___pip_5160_1_11___block_40_dt_y;
_q___pip_5160_1_12___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___block_40_dt_y : _d___pip_5160_1_12___block_40_dt_y;
_q___pip_5160_1_13___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___block_40_dt_y : _d___pip_5160_1_13___block_40_dt_y;
_q___pip_5160_1_14___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___block_40_dt_y : _d___pip_5160_1_14___block_40_dt_y;
_q___pip_5160_1_15___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___block_40_dt_y : _d___pip_5160_1_15___block_40_dt_y;
_q___pip_5160_1_16___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___block_40_dt_y : _d___pip_5160_1_16___block_40_dt_y;
_q___pip_5160_1_17___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___block_40_dt_y : _d___pip_5160_1_17___block_40_dt_y;
_q___pip_5160_1_18___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___block_40_dt_y : _d___pip_5160_1_18___block_40_dt_y;
_q___pip_5160_1_19___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___block_40_dt_y : _d___pip_5160_1_19___block_40_dt_y;
_q___pip_5160_1_20___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___block_40_dt_y : _d___pip_5160_1_20___block_40_dt_y;
_q___pip_5160_1_21___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___block_40_dt_y : _d___pip_5160_1_21___block_40_dt_y;
_q___pip_5160_1_22___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___block_40_dt_y : _d___pip_5160_1_22___block_40_dt_y;
_q___pip_5160_1_23___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___block_40_dt_y : _d___pip_5160_1_23___block_40_dt_y;
_q___pip_5160_1_24___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___block_40_dt_y : _d___pip_5160_1_24___block_40_dt_y;
_q___pip_5160_1_25___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___block_40_dt_y : _d___pip_5160_1_25___block_40_dt_y;
_q___pip_5160_1_26___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___block_40_dt_y : _d___pip_5160_1_26___block_40_dt_y;
_q___pip_5160_1_27___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___block_40_dt_y : _d___pip_5160_1_27___block_40_dt_y;
_q___pip_5160_1_28___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___block_40_dt_y : _d___pip_5160_1_28___block_40_dt_y;
_q___pip_5160_1_29___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___block_40_dt_y : _d___pip_5160_1_29___block_40_dt_y;
_q___pip_5160_1_30___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___block_40_dt_y : _d___pip_5160_1_30___block_40_dt_y;
_q___pip_5160_1_31___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___block_40_dt_y : _d___pip_5160_1_31___block_40_dt_y;
_q___pip_5160_1_32___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___block_40_dt_y : _d___pip_5160_1_32___block_40_dt_y;
_q___pip_5160_1_33___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___block_40_dt_y : _d___pip_5160_1_33___block_40_dt_y;
_q___pip_5160_1_34___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___block_40_dt_y : _d___pip_5160_1_34___block_40_dt_y;
_q___pip_5160_1_35___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___block_40_dt_y : _d___pip_5160_1_35___block_40_dt_y;
_q___pip_5160_1_36___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___block_40_dt_y : _d___pip_5160_1_36___block_40_dt_y;
_q___pip_5160_1_37___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___block_40_dt_y : _d___pip_5160_1_37___block_40_dt_y;
_q___pip_5160_1_38___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___block_40_dt_y : _d___pip_5160_1_38___block_40_dt_y;
_q___pip_5160_1_39___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___block_40_dt_y : _d___pip_5160_1_39___block_40_dt_y;
_q___pip_5160_1_40___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___block_40_dt_y : _d___pip_5160_1_40___block_40_dt_y;
_q___pip_5160_1_41___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___block_40_dt_y : _d___pip_5160_1_41___block_40_dt_y;
_q___pip_5160_1_42___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___block_40_dt_y : _d___pip_5160_1_42___block_40_dt_y;
_q___pip_5160_1_43___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___block_40_dt_y : _d___pip_5160_1_43___block_40_dt_y;
_q___pip_5160_1_44___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___block_40_dt_y : _d___pip_5160_1_44___block_40_dt_y;
_q___pip_5160_1_45___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___block_40_dt_y : _d___pip_5160_1_45___block_40_dt_y;
_q___pip_5160_1_46___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___block_40_dt_y : _d___pip_5160_1_46___block_40_dt_y;
_q___pip_5160_1_47___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___block_40_dt_y : _d___pip_5160_1_47___block_40_dt_y;
_q___pip_5160_1_48___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___block_40_dt_y : _d___pip_5160_1_48___block_40_dt_y;
_q___pip_5160_1_49___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___block_40_dt_y : _d___pip_5160_1_49___block_40_dt_y;
_q___pip_5160_1_50___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___block_40_dt_y : _d___pip_5160_1_50___block_40_dt_y;
_q___pip_5160_1_51___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___block_40_dt_y : _d___pip_5160_1_51___block_40_dt_y;
_q___pip_5160_1_52___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___block_40_dt_y : _d___pip_5160_1_52___block_40_dt_y;
_q___pip_5160_1_53___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___block_40_dt_y : _d___pip_5160_1_53___block_40_dt_y;
_q___pip_5160_1_54___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___block_40_dt_y : _d___pip_5160_1_54___block_40_dt_y;
_q___pip_5160_1_55___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___block_40_dt_y : _d___pip_5160_1_55___block_40_dt_y;
_q___pip_5160_1_56___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___block_40_dt_y : _d___pip_5160_1_56___block_40_dt_y;
_q___pip_5160_1_57___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___block_40_dt_y : _d___pip_5160_1_57___block_40_dt_y;
_q___pip_5160_1_58___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___block_40_dt_y : _d___pip_5160_1_58___block_40_dt_y;
_q___pip_5160_1_59___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___block_40_dt_y : _d___pip_5160_1_59___block_40_dt_y;
_q___pip_5160_1_60___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___block_40_dt_y : _d___pip_5160_1_60___block_40_dt_y;
_q___pip_5160_1_61___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___block_40_dt_y : _d___pip_5160_1_61___block_40_dt_y;
_q___pip_5160_1_62___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___block_40_dt_y : _d___pip_5160_1_62___block_40_dt_y;
_q___pip_5160_1_63___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___block_40_dt_y : _d___pip_5160_1_63___block_40_dt_y;
_q___pip_5160_1_64___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___block_40_dt_y : _d___pip_5160_1_64___block_40_dt_y;
_q___pip_5160_1_65___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___block_40_dt_y : _d___pip_5160_1_65___block_40_dt_y;
_q___pip_5160_1_66___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___block_40_dt_y : _d___pip_5160_1_66___block_40_dt_y;
_q___pip_5160_1_67___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___block_40_dt_y : _d___pip_5160_1_67___block_40_dt_y;
_q___pip_5160_1_68___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___block_40_dt_y : _d___pip_5160_1_68___block_40_dt_y;
_q___pip_5160_1_69___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___block_40_dt_y : _d___pip_5160_1_69___block_40_dt_y;
_q___pip_5160_1_70___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___block_40_dt_y : _d___pip_5160_1_70___block_40_dt_y;
_q___pip_5160_1_71___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___block_40_dt_y : _d___pip_5160_1_71___block_40_dt_y;
_q___pip_5160_1_72___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___block_40_dt_y : _d___pip_5160_1_72___block_40_dt_y;
_q___pip_5160_1_73___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___block_40_dt_y : _d___pip_5160_1_73___block_40_dt_y;
_q___pip_5160_1_74___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___block_40_dt_y : _d___pip_5160_1_74___block_40_dt_y;
_q___pip_5160_1_75___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___block_40_dt_y : _d___pip_5160_1_75___block_40_dt_y;
_q___pip_5160_1_76___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___block_40_dt_y : _d___pip_5160_1_76___block_40_dt_y;
_q___pip_5160_1_77___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___block_40_dt_y : _d___pip_5160_1_77___block_40_dt_y;
_q___pip_5160_1_78___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___block_40_dt_y : _d___pip_5160_1_78___block_40_dt_y;
_q___pip_5160_1_79___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___block_40_dt_y : _d___pip_5160_1_79___block_40_dt_y;
_q___pip_5160_1_80___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___block_40_dt_y : _d___pip_5160_1_80___block_40_dt_y;
_q___pip_5160_1_81___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___block_40_dt_y : _d___pip_5160_1_81___block_40_dt_y;
_q___pip_5160_1_82___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___block_40_dt_y : _d___pip_5160_1_82___block_40_dt_y;
_q___pip_5160_1_83___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___block_40_dt_y : _d___pip_5160_1_83___block_40_dt_y;
_q___pip_5160_1_84___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___block_40_dt_y : _d___pip_5160_1_84___block_40_dt_y;
_q___pip_5160_1_85___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___block_40_dt_y : _d___pip_5160_1_85___block_40_dt_y;
_q___pip_5160_1_86___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___block_40_dt_y : _d___pip_5160_1_86___block_40_dt_y;
_q___pip_5160_1_87___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___block_40_dt_y : _d___pip_5160_1_87___block_40_dt_y;
_q___pip_5160_1_88___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___block_40_dt_y : _d___pip_5160_1_88___block_40_dt_y;
_q___pip_5160_1_89___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___block_40_dt_y : _d___pip_5160_1_89___block_40_dt_y;
_q___pip_5160_1_90___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___block_40_dt_y : _d___pip_5160_1_90___block_40_dt_y;
_q___pip_5160_1_91___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___block_40_dt_y : _d___pip_5160_1_91___block_40_dt_y;
_q___pip_5160_1_92___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___block_40_dt_y : _d___pip_5160_1_92___block_40_dt_y;
_q___pip_5160_1_93___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___block_40_dt_y : _d___pip_5160_1_93___block_40_dt_y;
_q___pip_5160_1_94___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___block_40_dt_y : _d___pip_5160_1_94___block_40_dt_y;
_q___pip_5160_1_95___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___block_40_dt_y : _d___pip_5160_1_95___block_40_dt_y;
_q___pip_5160_1_96___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___block_40_dt_y : _d___pip_5160_1_96___block_40_dt_y;
_q___pip_5160_1_97___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___block_40_dt_y : _d___pip_5160_1_97___block_40_dt_y;
_q___pip_5160_1_98___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___block_40_dt_y : _d___pip_5160_1_98___block_40_dt_y;
_q___pip_5160_1_99___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___block_40_dt_y : _d___pip_5160_1_99___block_40_dt_y;
_q___pip_5160_1_100___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___block_40_dt_y : _d___pip_5160_1_100___block_40_dt_y;
_q___pip_5160_1_101___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___block_40_dt_y : _d___pip_5160_1_101___block_40_dt_y;
_q___pip_5160_1_102___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___block_40_dt_y : _d___pip_5160_1_102___block_40_dt_y;
_q___pip_5160_1_103___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___block_40_dt_y : _d___pip_5160_1_103___block_40_dt_y;
_q___pip_5160_1_104___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___block_40_dt_y : _d___pip_5160_1_104___block_40_dt_y;
_q___pip_5160_1_105___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___block_40_dt_y : _d___pip_5160_1_105___block_40_dt_y;
_q___pip_5160_1_106___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___block_40_dt_y : _d___pip_5160_1_106___block_40_dt_y;
_q___pip_5160_1_107___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___block_40_dt_y : _d___pip_5160_1_107___block_40_dt_y;
_q___pip_5160_1_108___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___block_40_dt_y : _d___pip_5160_1_108___block_40_dt_y;
_q___pip_5160_1_109___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___block_40_dt_y : _d___pip_5160_1_109___block_40_dt_y;
_q___pip_5160_1_110___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___block_40_dt_y : _d___pip_5160_1_110___block_40_dt_y;
_q___pip_5160_1_111___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___block_40_dt_y : _d___pip_5160_1_111___block_40_dt_y;
_q___pip_5160_1_112___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___block_40_dt_y : _d___pip_5160_1_112___block_40_dt_y;
_q___pip_5160_1_113___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___block_40_dt_y : _d___pip_5160_1_113___block_40_dt_y;
_q___pip_5160_1_114___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___block_40_dt_y : _d___pip_5160_1_114___block_40_dt_y;
_q___pip_5160_1_115___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___block_40_dt_y : _d___pip_5160_1_115___block_40_dt_y;
_q___pip_5160_1_116___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___block_40_dt_y : _d___pip_5160_1_116___block_40_dt_y;
_q___pip_5160_1_117___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___block_40_dt_y : _d___pip_5160_1_117___block_40_dt_y;
_q___pip_5160_1_118___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___block_40_dt_y : _d___pip_5160_1_118___block_40_dt_y;
_q___pip_5160_1_119___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___block_40_dt_y : _d___pip_5160_1_119___block_40_dt_y;
_q___pip_5160_1_120___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___block_40_dt_y : _d___pip_5160_1_120___block_40_dt_y;
_q___pip_5160_1_121___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___block_40_dt_y : _d___pip_5160_1_121___block_40_dt_y;
_q___pip_5160_1_122___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___block_40_dt_y : _d___pip_5160_1_122___block_40_dt_y;
_q___pip_5160_1_123___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___block_40_dt_y : _d___pip_5160_1_123___block_40_dt_y;
_q___pip_5160_1_124___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___block_40_dt_y : _d___pip_5160_1_124___block_40_dt_y;
_q___pip_5160_1_125___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___block_40_dt_y : _d___pip_5160_1_125___block_40_dt_y;
_q___pip_5160_1_126___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___block_40_dt_y : _d___pip_5160_1_126___block_40_dt_y;
_q___pip_5160_1_127___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___block_40_dt_y : _d___pip_5160_1_127___block_40_dt_y;
_q___pip_5160_1_128___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___block_40_dt_y : _d___pip_5160_1_128___block_40_dt_y;
_q___pip_5160_1_129___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___block_40_dt_y : _d___pip_5160_1_129___block_40_dt_y;
_q___pip_5160_1_130___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___block_40_dt_y : _d___pip_5160_1_130___block_40_dt_y;
_q___pip_5160_1_131___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___block_40_dt_y : _d___pip_5160_1_131___block_40_dt_y;
_q___pip_5160_1_132___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___block_40_dt_y : _d___pip_5160_1_132___block_40_dt_y;
_q___pip_5160_1_133___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___block_40_dt_y : _d___pip_5160_1_133___block_40_dt_y;
_q___pip_5160_1_134___block_40_dt_y <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___block_40_dt_y : _d___pip_5160_1_134___block_40_dt_y;
_q___pip_5160_1_6___block_40_dt_z <= _d___pip_5160_1_6___block_40_dt_z;
_q___pip_5160_1_7___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___block_40_dt_z : _d___pip_5160_1_7___block_40_dt_z;
_q___pip_5160_1_8___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___block_40_dt_z : _d___pip_5160_1_8___block_40_dt_z;
_q___pip_5160_1_9___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___block_40_dt_z : _d___pip_5160_1_9___block_40_dt_z;
_q___pip_5160_1_10___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___block_40_dt_z : _d___pip_5160_1_10___block_40_dt_z;
_q___pip_5160_1_11___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___block_40_dt_z : _d___pip_5160_1_11___block_40_dt_z;
_q___pip_5160_1_12___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___block_40_dt_z : _d___pip_5160_1_12___block_40_dt_z;
_q___pip_5160_1_13___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___block_40_dt_z : _d___pip_5160_1_13___block_40_dt_z;
_q___pip_5160_1_14___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___block_40_dt_z : _d___pip_5160_1_14___block_40_dt_z;
_q___pip_5160_1_15___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___block_40_dt_z : _d___pip_5160_1_15___block_40_dt_z;
_q___pip_5160_1_16___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___block_40_dt_z : _d___pip_5160_1_16___block_40_dt_z;
_q___pip_5160_1_17___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___block_40_dt_z : _d___pip_5160_1_17___block_40_dt_z;
_q___pip_5160_1_18___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___block_40_dt_z : _d___pip_5160_1_18___block_40_dt_z;
_q___pip_5160_1_19___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___block_40_dt_z : _d___pip_5160_1_19___block_40_dt_z;
_q___pip_5160_1_20___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___block_40_dt_z : _d___pip_5160_1_20___block_40_dt_z;
_q___pip_5160_1_21___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___block_40_dt_z : _d___pip_5160_1_21___block_40_dt_z;
_q___pip_5160_1_22___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___block_40_dt_z : _d___pip_5160_1_22___block_40_dt_z;
_q___pip_5160_1_23___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___block_40_dt_z : _d___pip_5160_1_23___block_40_dt_z;
_q___pip_5160_1_24___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___block_40_dt_z : _d___pip_5160_1_24___block_40_dt_z;
_q___pip_5160_1_25___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___block_40_dt_z : _d___pip_5160_1_25___block_40_dt_z;
_q___pip_5160_1_26___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___block_40_dt_z : _d___pip_5160_1_26___block_40_dt_z;
_q___pip_5160_1_27___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___block_40_dt_z : _d___pip_5160_1_27___block_40_dt_z;
_q___pip_5160_1_28___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___block_40_dt_z : _d___pip_5160_1_28___block_40_dt_z;
_q___pip_5160_1_29___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___block_40_dt_z : _d___pip_5160_1_29___block_40_dt_z;
_q___pip_5160_1_30___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___block_40_dt_z : _d___pip_5160_1_30___block_40_dt_z;
_q___pip_5160_1_31___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___block_40_dt_z : _d___pip_5160_1_31___block_40_dt_z;
_q___pip_5160_1_32___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___block_40_dt_z : _d___pip_5160_1_32___block_40_dt_z;
_q___pip_5160_1_33___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___block_40_dt_z : _d___pip_5160_1_33___block_40_dt_z;
_q___pip_5160_1_34___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___block_40_dt_z : _d___pip_5160_1_34___block_40_dt_z;
_q___pip_5160_1_35___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___block_40_dt_z : _d___pip_5160_1_35___block_40_dt_z;
_q___pip_5160_1_36___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___block_40_dt_z : _d___pip_5160_1_36___block_40_dt_z;
_q___pip_5160_1_37___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___block_40_dt_z : _d___pip_5160_1_37___block_40_dt_z;
_q___pip_5160_1_38___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___block_40_dt_z : _d___pip_5160_1_38___block_40_dt_z;
_q___pip_5160_1_39___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___block_40_dt_z : _d___pip_5160_1_39___block_40_dt_z;
_q___pip_5160_1_40___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___block_40_dt_z : _d___pip_5160_1_40___block_40_dt_z;
_q___pip_5160_1_41___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___block_40_dt_z : _d___pip_5160_1_41___block_40_dt_z;
_q___pip_5160_1_42___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___block_40_dt_z : _d___pip_5160_1_42___block_40_dt_z;
_q___pip_5160_1_43___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___block_40_dt_z : _d___pip_5160_1_43___block_40_dt_z;
_q___pip_5160_1_44___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___block_40_dt_z : _d___pip_5160_1_44___block_40_dt_z;
_q___pip_5160_1_45___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___block_40_dt_z : _d___pip_5160_1_45___block_40_dt_z;
_q___pip_5160_1_46___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___block_40_dt_z : _d___pip_5160_1_46___block_40_dt_z;
_q___pip_5160_1_47___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___block_40_dt_z : _d___pip_5160_1_47___block_40_dt_z;
_q___pip_5160_1_48___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___block_40_dt_z : _d___pip_5160_1_48___block_40_dt_z;
_q___pip_5160_1_49___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___block_40_dt_z : _d___pip_5160_1_49___block_40_dt_z;
_q___pip_5160_1_50___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___block_40_dt_z : _d___pip_5160_1_50___block_40_dt_z;
_q___pip_5160_1_51___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___block_40_dt_z : _d___pip_5160_1_51___block_40_dt_z;
_q___pip_5160_1_52___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___block_40_dt_z : _d___pip_5160_1_52___block_40_dt_z;
_q___pip_5160_1_53___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___block_40_dt_z : _d___pip_5160_1_53___block_40_dt_z;
_q___pip_5160_1_54___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___block_40_dt_z : _d___pip_5160_1_54___block_40_dt_z;
_q___pip_5160_1_55___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___block_40_dt_z : _d___pip_5160_1_55___block_40_dt_z;
_q___pip_5160_1_56___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___block_40_dt_z : _d___pip_5160_1_56___block_40_dt_z;
_q___pip_5160_1_57___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___block_40_dt_z : _d___pip_5160_1_57___block_40_dt_z;
_q___pip_5160_1_58___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___block_40_dt_z : _d___pip_5160_1_58___block_40_dt_z;
_q___pip_5160_1_59___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___block_40_dt_z : _d___pip_5160_1_59___block_40_dt_z;
_q___pip_5160_1_60___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___block_40_dt_z : _d___pip_5160_1_60___block_40_dt_z;
_q___pip_5160_1_61___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___block_40_dt_z : _d___pip_5160_1_61___block_40_dt_z;
_q___pip_5160_1_62___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___block_40_dt_z : _d___pip_5160_1_62___block_40_dt_z;
_q___pip_5160_1_63___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___block_40_dt_z : _d___pip_5160_1_63___block_40_dt_z;
_q___pip_5160_1_64___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___block_40_dt_z : _d___pip_5160_1_64___block_40_dt_z;
_q___pip_5160_1_65___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___block_40_dt_z : _d___pip_5160_1_65___block_40_dt_z;
_q___pip_5160_1_66___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___block_40_dt_z : _d___pip_5160_1_66___block_40_dt_z;
_q___pip_5160_1_67___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___block_40_dt_z : _d___pip_5160_1_67___block_40_dt_z;
_q___pip_5160_1_68___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___block_40_dt_z : _d___pip_5160_1_68___block_40_dt_z;
_q___pip_5160_1_69___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___block_40_dt_z : _d___pip_5160_1_69___block_40_dt_z;
_q___pip_5160_1_70___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___block_40_dt_z : _d___pip_5160_1_70___block_40_dt_z;
_q___pip_5160_1_71___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___block_40_dt_z : _d___pip_5160_1_71___block_40_dt_z;
_q___pip_5160_1_72___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___block_40_dt_z : _d___pip_5160_1_72___block_40_dt_z;
_q___pip_5160_1_73___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___block_40_dt_z : _d___pip_5160_1_73___block_40_dt_z;
_q___pip_5160_1_74___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___block_40_dt_z : _d___pip_5160_1_74___block_40_dt_z;
_q___pip_5160_1_75___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___block_40_dt_z : _d___pip_5160_1_75___block_40_dt_z;
_q___pip_5160_1_76___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___block_40_dt_z : _d___pip_5160_1_76___block_40_dt_z;
_q___pip_5160_1_77___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___block_40_dt_z : _d___pip_5160_1_77___block_40_dt_z;
_q___pip_5160_1_78___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___block_40_dt_z : _d___pip_5160_1_78___block_40_dt_z;
_q___pip_5160_1_79___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___block_40_dt_z : _d___pip_5160_1_79___block_40_dt_z;
_q___pip_5160_1_80___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___block_40_dt_z : _d___pip_5160_1_80___block_40_dt_z;
_q___pip_5160_1_81___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___block_40_dt_z : _d___pip_5160_1_81___block_40_dt_z;
_q___pip_5160_1_82___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___block_40_dt_z : _d___pip_5160_1_82___block_40_dt_z;
_q___pip_5160_1_83___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___block_40_dt_z : _d___pip_5160_1_83___block_40_dt_z;
_q___pip_5160_1_84___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___block_40_dt_z : _d___pip_5160_1_84___block_40_dt_z;
_q___pip_5160_1_85___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___block_40_dt_z : _d___pip_5160_1_85___block_40_dt_z;
_q___pip_5160_1_86___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___block_40_dt_z : _d___pip_5160_1_86___block_40_dt_z;
_q___pip_5160_1_87___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___block_40_dt_z : _d___pip_5160_1_87___block_40_dt_z;
_q___pip_5160_1_88___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___block_40_dt_z : _d___pip_5160_1_88___block_40_dt_z;
_q___pip_5160_1_89___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___block_40_dt_z : _d___pip_5160_1_89___block_40_dt_z;
_q___pip_5160_1_90___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___block_40_dt_z : _d___pip_5160_1_90___block_40_dt_z;
_q___pip_5160_1_91___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___block_40_dt_z : _d___pip_5160_1_91___block_40_dt_z;
_q___pip_5160_1_92___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___block_40_dt_z : _d___pip_5160_1_92___block_40_dt_z;
_q___pip_5160_1_93___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___block_40_dt_z : _d___pip_5160_1_93___block_40_dt_z;
_q___pip_5160_1_94___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___block_40_dt_z : _d___pip_5160_1_94___block_40_dt_z;
_q___pip_5160_1_95___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___block_40_dt_z : _d___pip_5160_1_95___block_40_dt_z;
_q___pip_5160_1_96___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___block_40_dt_z : _d___pip_5160_1_96___block_40_dt_z;
_q___pip_5160_1_97___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___block_40_dt_z : _d___pip_5160_1_97___block_40_dt_z;
_q___pip_5160_1_98___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___block_40_dt_z : _d___pip_5160_1_98___block_40_dt_z;
_q___pip_5160_1_99___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___block_40_dt_z : _d___pip_5160_1_99___block_40_dt_z;
_q___pip_5160_1_100___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___block_40_dt_z : _d___pip_5160_1_100___block_40_dt_z;
_q___pip_5160_1_101___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___block_40_dt_z : _d___pip_5160_1_101___block_40_dt_z;
_q___pip_5160_1_102___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___block_40_dt_z : _d___pip_5160_1_102___block_40_dt_z;
_q___pip_5160_1_103___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___block_40_dt_z : _d___pip_5160_1_103___block_40_dt_z;
_q___pip_5160_1_104___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___block_40_dt_z : _d___pip_5160_1_104___block_40_dt_z;
_q___pip_5160_1_105___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___block_40_dt_z : _d___pip_5160_1_105___block_40_dt_z;
_q___pip_5160_1_106___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___block_40_dt_z : _d___pip_5160_1_106___block_40_dt_z;
_q___pip_5160_1_107___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___block_40_dt_z : _d___pip_5160_1_107___block_40_dt_z;
_q___pip_5160_1_108___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___block_40_dt_z : _d___pip_5160_1_108___block_40_dt_z;
_q___pip_5160_1_109___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___block_40_dt_z : _d___pip_5160_1_109___block_40_dt_z;
_q___pip_5160_1_110___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___block_40_dt_z : _d___pip_5160_1_110___block_40_dt_z;
_q___pip_5160_1_111___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___block_40_dt_z : _d___pip_5160_1_111___block_40_dt_z;
_q___pip_5160_1_112___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___block_40_dt_z : _d___pip_5160_1_112___block_40_dt_z;
_q___pip_5160_1_113___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___block_40_dt_z : _d___pip_5160_1_113___block_40_dt_z;
_q___pip_5160_1_114___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___block_40_dt_z : _d___pip_5160_1_114___block_40_dt_z;
_q___pip_5160_1_115___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___block_40_dt_z : _d___pip_5160_1_115___block_40_dt_z;
_q___pip_5160_1_116___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___block_40_dt_z : _d___pip_5160_1_116___block_40_dt_z;
_q___pip_5160_1_117___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___block_40_dt_z : _d___pip_5160_1_117___block_40_dt_z;
_q___pip_5160_1_118___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___block_40_dt_z : _d___pip_5160_1_118___block_40_dt_z;
_q___pip_5160_1_119___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___block_40_dt_z : _d___pip_5160_1_119___block_40_dt_z;
_q___pip_5160_1_120___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___block_40_dt_z : _d___pip_5160_1_120___block_40_dt_z;
_q___pip_5160_1_121___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___block_40_dt_z : _d___pip_5160_1_121___block_40_dt_z;
_q___pip_5160_1_122___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___block_40_dt_z : _d___pip_5160_1_122___block_40_dt_z;
_q___pip_5160_1_123___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___block_40_dt_z : _d___pip_5160_1_123___block_40_dt_z;
_q___pip_5160_1_124___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___block_40_dt_z : _d___pip_5160_1_124___block_40_dt_z;
_q___pip_5160_1_125___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___block_40_dt_z : _d___pip_5160_1_125___block_40_dt_z;
_q___pip_5160_1_126___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___block_40_dt_z : _d___pip_5160_1_126___block_40_dt_z;
_q___pip_5160_1_127___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___block_40_dt_z : _d___pip_5160_1_127___block_40_dt_z;
_q___pip_5160_1_128___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___block_40_dt_z : _d___pip_5160_1_128___block_40_dt_z;
_q___pip_5160_1_129___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___block_40_dt_z : _d___pip_5160_1_129___block_40_dt_z;
_q___pip_5160_1_130___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___block_40_dt_z : _d___pip_5160_1_130___block_40_dt_z;
_q___pip_5160_1_131___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___block_40_dt_z : _d___pip_5160_1_131___block_40_dt_z;
_q___pip_5160_1_132___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___block_40_dt_z : _d___pip_5160_1_132___block_40_dt_z;
_q___pip_5160_1_133___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___block_40_dt_z : _d___pip_5160_1_133___block_40_dt_z;
_q___pip_5160_1_134___block_40_dt_z <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___block_40_dt_z : _d___pip_5160_1_134___block_40_dt_z;
_q___pip_5160_1_4___stage___block_26_brd_x <= _d___pip_5160_1_4___stage___block_26_brd_x;
_q___pip_5160_1_5___stage___block_26_brd_x <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_26_brd_x : _d___pip_5160_1_5___stage___block_26_brd_x;
_q___pip_5160_1_6___stage___block_26_brd_x <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_26_brd_x : _d___pip_5160_1_6___stage___block_26_brd_x;
_q___pip_5160_1_4___stage___block_26_brd_y <= _d___pip_5160_1_4___stage___block_26_brd_y;
_q___pip_5160_1_5___stage___block_26_brd_y <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_26_brd_y : _d___pip_5160_1_5___stage___block_26_brd_y;
_q___pip_5160_1_6___stage___block_26_brd_y <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_26_brd_y : _d___pip_5160_1_6___stage___block_26_brd_y;
_q___pip_5160_1_4___stage___block_26_brd_z <= _d___pip_5160_1_4___stage___block_26_brd_z;
_q___pip_5160_1_5___stage___block_26_brd_z <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_26_brd_z : _d___pip_5160_1_5___stage___block_26_brd_z;
_q___pip_5160_1_6___stage___block_26_brd_z <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_26_brd_z : _d___pip_5160_1_6___stage___block_26_brd_z;
_q___pip_5160_1_4___stage___block_26_rd_x <= _d___pip_5160_1_4___stage___block_26_rd_x;
_q___pip_5160_1_5___stage___block_26_rd_x <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_26_rd_x : _d___pip_5160_1_5___stage___block_26_rd_x;
_q___pip_5160_1_4___stage___block_26_rd_y <= _d___pip_5160_1_4___stage___block_26_rd_y;
_q___pip_5160_1_5___stage___block_26_rd_y <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_26_rd_y : _d___pip_5160_1_5___stage___block_26_rd_y;
_q___pip_5160_1_4___stage___block_26_rd_z <= _d___pip_5160_1_4___stage___block_26_rd_z;
_q___pip_5160_1_5___stage___block_26_rd_z <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_26_rd_z : _d___pip_5160_1_5___stage___block_26_rd_z;
_q___pip_5160_1_4___stage___block_26_s_x <= _d___pip_5160_1_4___stage___block_26_s_x;
_q___pip_5160_1_5___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_26_s_x : _d___pip_5160_1_5___stage___block_26_s_x;
_q___pip_5160_1_6___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_26_s_x : _d___pip_5160_1_6___stage___block_26_s_x;
_q___pip_5160_1_7___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___stage___block_26_s_x : _d___pip_5160_1_7___stage___block_26_s_x;
_q___pip_5160_1_8___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___stage___block_26_s_x : _d___pip_5160_1_8___stage___block_26_s_x;
_q___pip_5160_1_9___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___stage___block_26_s_x : _d___pip_5160_1_9___stage___block_26_s_x;
_q___pip_5160_1_10___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___stage___block_26_s_x : _d___pip_5160_1_10___stage___block_26_s_x;
_q___pip_5160_1_11___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___stage___block_26_s_x : _d___pip_5160_1_11___stage___block_26_s_x;
_q___pip_5160_1_12___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___stage___block_26_s_x : _d___pip_5160_1_12___stage___block_26_s_x;
_q___pip_5160_1_13___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___stage___block_26_s_x : _d___pip_5160_1_13___stage___block_26_s_x;
_q___pip_5160_1_14___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___stage___block_26_s_x : _d___pip_5160_1_14___stage___block_26_s_x;
_q___pip_5160_1_15___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___stage___block_26_s_x : _d___pip_5160_1_15___stage___block_26_s_x;
_q___pip_5160_1_16___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___stage___block_26_s_x : _d___pip_5160_1_16___stage___block_26_s_x;
_q___pip_5160_1_17___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___stage___block_26_s_x : _d___pip_5160_1_17___stage___block_26_s_x;
_q___pip_5160_1_18___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___stage___block_26_s_x : _d___pip_5160_1_18___stage___block_26_s_x;
_q___pip_5160_1_19___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___stage___block_26_s_x : _d___pip_5160_1_19___stage___block_26_s_x;
_q___pip_5160_1_20___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___stage___block_26_s_x : _d___pip_5160_1_20___stage___block_26_s_x;
_q___pip_5160_1_21___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___stage___block_26_s_x : _d___pip_5160_1_21___stage___block_26_s_x;
_q___pip_5160_1_22___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___stage___block_26_s_x : _d___pip_5160_1_22___stage___block_26_s_x;
_q___pip_5160_1_23___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___stage___block_26_s_x : _d___pip_5160_1_23___stage___block_26_s_x;
_q___pip_5160_1_24___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___stage___block_26_s_x : _d___pip_5160_1_24___stage___block_26_s_x;
_q___pip_5160_1_25___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___stage___block_26_s_x : _d___pip_5160_1_25___stage___block_26_s_x;
_q___pip_5160_1_26___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___stage___block_26_s_x : _d___pip_5160_1_26___stage___block_26_s_x;
_q___pip_5160_1_27___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___stage___block_26_s_x : _d___pip_5160_1_27___stage___block_26_s_x;
_q___pip_5160_1_28___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___stage___block_26_s_x : _d___pip_5160_1_28___stage___block_26_s_x;
_q___pip_5160_1_29___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___stage___block_26_s_x : _d___pip_5160_1_29___stage___block_26_s_x;
_q___pip_5160_1_30___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___stage___block_26_s_x : _d___pip_5160_1_30___stage___block_26_s_x;
_q___pip_5160_1_31___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___stage___block_26_s_x : _d___pip_5160_1_31___stage___block_26_s_x;
_q___pip_5160_1_32___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___stage___block_26_s_x : _d___pip_5160_1_32___stage___block_26_s_x;
_q___pip_5160_1_33___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___stage___block_26_s_x : _d___pip_5160_1_33___stage___block_26_s_x;
_q___pip_5160_1_34___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___stage___block_26_s_x : _d___pip_5160_1_34___stage___block_26_s_x;
_q___pip_5160_1_35___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___stage___block_26_s_x : _d___pip_5160_1_35___stage___block_26_s_x;
_q___pip_5160_1_36___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___stage___block_26_s_x : _d___pip_5160_1_36___stage___block_26_s_x;
_q___pip_5160_1_37___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___stage___block_26_s_x : _d___pip_5160_1_37___stage___block_26_s_x;
_q___pip_5160_1_38___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___stage___block_26_s_x : _d___pip_5160_1_38___stage___block_26_s_x;
_q___pip_5160_1_39___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___stage___block_26_s_x : _d___pip_5160_1_39___stage___block_26_s_x;
_q___pip_5160_1_40___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___stage___block_26_s_x : _d___pip_5160_1_40___stage___block_26_s_x;
_q___pip_5160_1_41___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___stage___block_26_s_x : _d___pip_5160_1_41___stage___block_26_s_x;
_q___pip_5160_1_42___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___stage___block_26_s_x : _d___pip_5160_1_42___stage___block_26_s_x;
_q___pip_5160_1_43___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___stage___block_26_s_x : _d___pip_5160_1_43___stage___block_26_s_x;
_q___pip_5160_1_44___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___stage___block_26_s_x : _d___pip_5160_1_44___stage___block_26_s_x;
_q___pip_5160_1_45___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___stage___block_26_s_x : _d___pip_5160_1_45___stage___block_26_s_x;
_q___pip_5160_1_46___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___stage___block_26_s_x : _d___pip_5160_1_46___stage___block_26_s_x;
_q___pip_5160_1_47___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___stage___block_26_s_x : _d___pip_5160_1_47___stage___block_26_s_x;
_q___pip_5160_1_48___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___stage___block_26_s_x : _d___pip_5160_1_48___stage___block_26_s_x;
_q___pip_5160_1_49___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___stage___block_26_s_x : _d___pip_5160_1_49___stage___block_26_s_x;
_q___pip_5160_1_50___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___stage___block_26_s_x : _d___pip_5160_1_50___stage___block_26_s_x;
_q___pip_5160_1_51___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___stage___block_26_s_x : _d___pip_5160_1_51___stage___block_26_s_x;
_q___pip_5160_1_52___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___stage___block_26_s_x : _d___pip_5160_1_52___stage___block_26_s_x;
_q___pip_5160_1_53___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___stage___block_26_s_x : _d___pip_5160_1_53___stage___block_26_s_x;
_q___pip_5160_1_54___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___stage___block_26_s_x : _d___pip_5160_1_54___stage___block_26_s_x;
_q___pip_5160_1_55___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___stage___block_26_s_x : _d___pip_5160_1_55___stage___block_26_s_x;
_q___pip_5160_1_56___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___stage___block_26_s_x : _d___pip_5160_1_56___stage___block_26_s_x;
_q___pip_5160_1_57___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___stage___block_26_s_x : _d___pip_5160_1_57___stage___block_26_s_x;
_q___pip_5160_1_58___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___stage___block_26_s_x : _d___pip_5160_1_58___stage___block_26_s_x;
_q___pip_5160_1_59___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___stage___block_26_s_x : _d___pip_5160_1_59___stage___block_26_s_x;
_q___pip_5160_1_60___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___stage___block_26_s_x : _d___pip_5160_1_60___stage___block_26_s_x;
_q___pip_5160_1_61___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___stage___block_26_s_x : _d___pip_5160_1_61___stage___block_26_s_x;
_q___pip_5160_1_62___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___stage___block_26_s_x : _d___pip_5160_1_62___stage___block_26_s_x;
_q___pip_5160_1_63___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___stage___block_26_s_x : _d___pip_5160_1_63___stage___block_26_s_x;
_q___pip_5160_1_64___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___stage___block_26_s_x : _d___pip_5160_1_64___stage___block_26_s_x;
_q___pip_5160_1_65___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___stage___block_26_s_x : _d___pip_5160_1_65___stage___block_26_s_x;
_q___pip_5160_1_66___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___stage___block_26_s_x : _d___pip_5160_1_66___stage___block_26_s_x;
_q___pip_5160_1_67___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___stage___block_26_s_x : _d___pip_5160_1_67___stage___block_26_s_x;
_q___pip_5160_1_68___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___stage___block_26_s_x : _d___pip_5160_1_68___stage___block_26_s_x;
_q___pip_5160_1_69___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___stage___block_26_s_x : _d___pip_5160_1_69___stage___block_26_s_x;
_q___pip_5160_1_70___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___stage___block_26_s_x : _d___pip_5160_1_70___stage___block_26_s_x;
_q___pip_5160_1_71___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___stage___block_26_s_x : _d___pip_5160_1_71___stage___block_26_s_x;
_q___pip_5160_1_72___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___stage___block_26_s_x : _d___pip_5160_1_72___stage___block_26_s_x;
_q___pip_5160_1_73___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___stage___block_26_s_x : _d___pip_5160_1_73___stage___block_26_s_x;
_q___pip_5160_1_74___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___stage___block_26_s_x : _d___pip_5160_1_74___stage___block_26_s_x;
_q___pip_5160_1_75___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___stage___block_26_s_x : _d___pip_5160_1_75___stage___block_26_s_x;
_q___pip_5160_1_76___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___stage___block_26_s_x : _d___pip_5160_1_76___stage___block_26_s_x;
_q___pip_5160_1_77___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___stage___block_26_s_x : _d___pip_5160_1_77___stage___block_26_s_x;
_q___pip_5160_1_78___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___stage___block_26_s_x : _d___pip_5160_1_78___stage___block_26_s_x;
_q___pip_5160_1_79___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___stage___block_26_s_x : _d___pip_5160_1_79___stage___block_26_s_x;
_q___pip_5160_1_80___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___stage___block_26_s_x : _d___pip_5160_1_80___stage___block_26_s_x;
_q___pip_5160_1_81___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___stage___block_26_s_x : _d___pip_5160_1_81___stage___block_26_s_x;
_q___pip_5160_1_82___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___stage___block_26_s_x : _d___pip_5160_1_82___stage___block_26_s_x;
_q___pip_5160_1_83___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___stage___block_26_s_x : _d___pip_5160_1_83___stage___block_26_s_x;
_q___pip_5160_1_84___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___stage___block_26_s_x : _d___pip_5160_1_84___stage___block_26_s_x;
_q___pip_5160_1_85___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___stage___block_26_s_x : _d___pip_5160_1_85___stage___block_26_s_x;
_q___pip_5160_1_86___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___stage___block_26_s_x : _d___pip_5160_1_86___stage___block_26_s_x;
_q___pip_5160_1_87___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___stage___block_26_s_x : _d___pip_5160_1_87___stage___block_26_s_x;
_q___pip_5160_1_88___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___stage___block_26_s_x : _d___pip_5160_1_88___stage___block_26_s_x;
_q___pip_5160_1_89___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___stage___block_26_s_x : _d___pip_5160_1_89___stage___block_26_s_x;
_q___pip_5160_1_90___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___stage___block_26_s_x : _d___pip_5160_1_90___stage___block_26_s_x;
_q___pip_5160_1_91___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___stage___block_26_s_x : _d___pip_5160_1_91___stage___block_26_s_x;
_q___pip_5160_1_92___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___stage___block_26_s_x : _d___pip_5160_1_92___stage___block_26_s_x;
_q___pip_5160_1_93___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___stage___block_26_s_x : _d___pip_5160_1_93___stage___block_26_s_x;
_q___pip_5160_1_94___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___stage___block_26_s_x : _d___pip_5160_1_94___stage___block_26_s_x;
_q___pip_5160_1_95___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___stage___block_26_s_x : _d___pip_5160_1_95___stage___block_26_s_x;
_q___pip_5160_1_96___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___stage___block_26_s_x : _d___pip_5160_1_96___stage___block_26_s_x;
_q___pip_5160_1_97___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___stage___block_26_s_x : _d___pip_5160_1_97___stage___block_26_s_x;
_q___pip_5160_1_98___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___stage___block_26_s_x : _d___pip_5160_1_98___stage___block_26_s_x;
_q___pip_5160_1_99___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___stage___block_26_s_x : _d___pip_5160_1_99___stage___block_26_s_x;
_q___pip_5160_1_100___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___stage___block_26_s_x : _d___pip_5160_1_100___stage___block_26_s_x;
_q___pip_5160_1_101___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___stage___block_26_s_x : _d___pip_5160_1_101___stage___block_26_s_x;
_q___pip_5160_1_102___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___stage___block_26_s_x : _d___pip_5160_1_102___stage___block_26_s_x;
_q___pip_5160_1_103___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___stage___block_26_s_x : _d___pip_5160_1_103___stage___block_26_s_x;
_q___pip_5160_1_104___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___stage___block_26_s_x : _d___pip_5160_1_104___stage___block_26_s_x;
_q___pip_5160_1_105___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___stage___block_26_s_x : _d___pip_5160_1_105___stage___block_26_s_x;
_q___pip_5160_1_106___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___stage___block_26_s_x : _d___pip_5160_1_106___stage___block_26_s_x;
_q___pip_5160_1_107___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___stage___block_26_s_x : _d___pip_5160_1_107___stage___block_26_s_x;
_q___pip_5160_1_108___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___stage___block_26_s_x : _d___pip_5160_1_108___stage___block_26_s_x;
_q___pip_5160_1_109___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___stage___block_26_s_x : _d___pip_5160_1_109___stage___block_26_s_x;
_q___pip_5160_1_110___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___stage___block_26_s_x : _d___pip_5160_1_110___stage___block_26_s_x;
_q___pip_5160_1_111___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___stage___block_26_s_x : _d___pip_5160_1_111___stage___block_26_s_x;
_q___pip_5160_1_112___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___stage___block_26_s_x : _d___pip_5160_1_112___stage___block_26_s_x;
_q___pip_5160_1_113___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___stage___block_26_s_x : _d___pip_5160_1_113___stage___block_26_s_x;
_q___pip_5160_1_114___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___stage___block_26_s_x : _d___pip_5160_1_114___stage___block_26_s_x;
_q___pip_5160_1_115___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___stage___block_26_s_x : _d___pip_5160_1_115___stage___block_26_s_x;
_q___pip_5160_1_116___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___stage___block_26_s_x : _d___pip_5160_1_116___stage___block_26_s_x;
_q___pip_5160_1_117___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___stage___block_26_s_x : _d___pip_5160_1_117___stage___block_26_s_x;
_q___pip_5160_1_118___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___stage___block_26_s_x : _d___pip_5160_1_118___stage___block_26_s_x;
_q___pip_5160_1_119___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___stage___block_26_s_x : _d___pip_5160_1_119___stage___block_26_s_x;
_q___pip_5160_1_120___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___stage___block_26_s_x : _d___pip_5160_1_120___stage___block_26_s_x;
_q___pip_5160_1_121___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___stage___block_26_s_x : _d___pip_5160_1_121___stage___block_26_s_x;
_q___pip_5160_1_122___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___stage___block_26_s_x : _d___pip_5160_1_122___stage___block_26_s_x;
_q___pip_5160_1_123___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___stage___block_26_s_x : _d___pip_5160_1_123___stage___block_26_s_x;
_q___pip_5160_1_124___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___stage___block_26_s_x : _d___pip_5160_1_124___stage___block_26_s_x;
_q___pip_5160_1_125___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___stage___block_26_s_x : _d___pip_5160_1_125___stage___block_26_s_x;
_q___pip_5160_1_126___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___stage___block_26_s_x : _d___pip_5160_1_126___stage___block_26_s_x;
_q___pip_5160_1_127___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___stage___block_26_s_x : _d___pip_5160_1_127___stage___block_26_s_x;
_q___pip_5160_1_128___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___stage___block_26_s_x : _d___pip_5160_1_128___stage___block_26_s_x;
_q___pip_5160_1_129___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___stage___block_26_s_x : _d___pip_5160_1_129___stage___block_26_s_x;
_q___pip_5160_1_130___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___stage___block_26_s_x : _d___pip_5160_1_130___stage___block_26_s_x;
_q___pip_5160_1_131___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___stage___block_26_s_x : _d___pip_5160_1_131___stage___block_26_s_x;
_q___pip_5160_1_132___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___stage___block_26_s_x : _d___pip_5160_1_132___stage___block_26_s_x;
_q___pip_5160_1_133___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___stage___block_26_s_x : _d___pip_5160_1_133___stage___block_26_s_x;
_q___pip_5160_1_134___stage___block_26_s_x <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___stage___block_26_s_x : _d___pip_5160_1_134___stage___block_26_s_x;
_q___pip_5160_1_4___stage___block_26_s_y <= _d___pip_5160_1_4___stage___block_26_s_y;
_q___pip_5160_1_5___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_26_s_y : _d___pip_5160_1_5___stage___block_26_s_y;
_q___pip_5160_1_6___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_26_s_y : _d___pip_5160_1_6___stage___block_26_s_y;
_q___pip_5160_1_7___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___stage___block_26_s_y : _d___pip_5160_1_7___stage___block_26_s_y;
_q___pip_5160_1_8___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___stage___block_26_s_y : _d___pip_5160_1_8___stage___block_26_s_y;
_q___pip_5160_1_9___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___stage___block_26_s_y : _d___pip_5160_1_9___stage___block_26_s_y;
_q___pip_5160_1_10___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___stage___block_26_s_y : _d___pip_5160_1_10___stage___block_26_s_y;
_q___pip_5160_1_11___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___stage___block_26_s_y : _d___pip_5160_1_11___stage___block_26_s_y;
_q___pip_5160_1_12___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___stage___block_26_s_y : _d___pip_5160_1_12___stage___block_26_s_y;
_q___pip_5160_1_13___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___stage___block_26_s_y : _d___pip_5160_1_13___stage___block_26_s_y;
_q___pip_5160_1_14___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___stage___block_26_s_y : _d___pip_5160_1_14___stage___block_26_s_y;
_q___pip_5160_1_15___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___stage___block_26_s_y : _d___pip_5160_1_15___stage___block_26_s_y;
_q___pip_5160_1_16___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___stage___block_26_s_y : _d___pip_5160_1_16___stage___block_26_s_y;
_q___pip_5160_1_17___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___stage___block_26_s_y : _d___pip_5160_1_17___stage___block_26_s_y;
_q___pip_5160_1_18___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___stage___block_26_s_y : _d___pip_5160_1_18___stage___block_26_s_y;
_q___pip_5160_1_19___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___stage___block_26_s_y : _d___pip_5160_1_19___stage___block_26_s_y;
_q___pip_5160_1_20___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___stage___block_26_s_y : _d___pip_5160_1_20___stage___block_26_s_y;
_q___pip_5160_1_21___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___stage___block_26_s_y : _d___pip_5160_1_21___stage___block_26_s_y;
_q___pip_5160_1_22___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___stage___block_26_s_y : _d___pip_5160_1_22___stage___block_26_s_y;
_q___pip_5160_1_23___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___stage___block_26_s_y : _d___pip_5160_1_23___stage___block_26_s_y;
_q___pip_5160_1_24___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___stage___block_26_s_y : _d___pip_5160_1_24___stage___block_26_s_y;
_q___pip_5160_1_25___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___stage___block_26_s_y : _d___pip_5160_1_25___stage___block_26_s_y;
_q___pip_5160_1_26___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___stage___block_26_s_y : _d___pip_5160_1_26___stage___block_26_s_y;
_q___pip_5160_1_27___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___stage___block_26_s_y : _d___pip_5160_1_27___stage___block_26_s_y;
_q___pip_5160_1_28___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___stage___block_26_s_y : _d___pip_5160_1_28___stage___block_26_s_y;
_q___pip_5160_1_29___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___stage___block_26_s_y : _d___pip_5160_1_29___stage___block_26_s_y;
_q___pip_5160_1_30___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___stage___block_26_s_y : _d___pip_5160_1_30___stage___block_26_s_y;
_q___pip_5160_1_31___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___stage___block_26_s_y : _d___pip_5160_1_31___stage___block_26_s_y;
_q___pip_5160_1_32___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___stage___block_26_s_y : _d___pip_5160_1_32___stage___block_26_s_y;
_q___pip_5160_1_33___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___stage___block_26_s_y : _d___pip_5160_1_33___stage___block_26_s_y;
_q___pip_5160_1_34___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___stage___block_26_s_y : _d___pip_5160_1_34___stage___block_26_s_y;
_q___pip_5160_1_35___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___stage___block_26_s_y : _d___pip_5160_1_35___stage___block_26_s_y;
_q___pip_5160_1_36___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___stage___block_26_s_y : _d___pip_5160_1_36___stage___block_26_s_y;
_q___pip_5160_1_37___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___stage___block_26_s_y : _d___pip_5160_1_37___stage___block_26_s_y;
_q___pip_5160_1_38___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___stage___block_26_s_y : _d___pip_5160_1_38___stage___block_26_s_y;
_q___pip_5160_1_39___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___stage___block_26_s_y : _d___pip_5160_1_39___stage___block_26_s_y;
_q___pip_5160_1_40___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___stage___block_26_s_y : _d___pip_5160_1_40___stage___block_26_s_y;
_q___pip_5160_1_41___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___stage___block_26_s_y : _d___pip_5160_1_41___stage___block_26_s_y;
_q___pip_5160_1_42___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___stage___block_26_s_y : _d___pip_5160_1_42___stage___block_26_s_y;
_q___pip_5160_1_43___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___stage___block_26_s_y : _d___pip_5160_1_43___stage___block_26_s_y;
_q___pip_5160_1_44___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___stage___block_26_s_y : _d___pip_5160_1_44___stage___block_26_s_y;
_q___pip_5160_1_45___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___stage___block_26_s_y : _d___pip_5160_1_45___stage___block_26_s_y;
_q___pip_5160_1_46___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___stage___block_26_s_y : _d___pip_5160_1_46___stage___block_26_s_y;
_q___pip_5160_1_47___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___stage___block_26_s_y : _d___pip_5160_1_47___stage___block_26_s_y;
_q___pip_5160_1_48___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___stage___block_26_s_y : _d___pip_5160_1_48___stage___block_26_s_y;
_q___pip_5160_1_49___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___stage___block_26_s_y : _d___pip_5160_1_49___stage___block_26_s_y;
_q___pip_5160_1_50___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___stage___block_26_s_y : _d___pip_5160_1_50___stage___block_26_s_y;
_q___pip_5160_1_51___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___stage___block_26_s_y : _d___pip_5160_1_51___stage___block_26_s_y;
_q___pip_5160_1_52___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___stage___block_26_s_y : _d___pip_5160_1_52___stage___block_26_s_y;
_q___pip_5160_1_53___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___stage___block_26_s_y : _d___pip_5160_1_53___stage___block_26_s_y;
_q___pip_5160_1_54___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___stage___block_26_s_y : _d___pip_5160_1_54___stage___block_26_s_y;
_q___pip_5160_1_55___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___stage___block_26_s_y : _d___pip_5160_1_55___stage___block_26_s_y;
_q___pip_5160_1_56___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___stage___block_26_s_y : _d___pip_5160_1_56___stage___block_26_s_y;
_q___pip_5160_1_57___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___stage___block_26_s_y : _d___pip_5160_1_57___stage___block_26_s_y;
_q___pip_5160_1_58___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___stage___block_26_s_y : _d___pip_5160_1_58___stage___block_26_s_y;
_q___pip_5160_1_59___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___stage___block_26_s_y : _d___pip_5160_1_59___stage___block_26_s_y;
_q___pip_5160_1_60___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___stage___block_26_s_y : _d___pip_5160_1_60___stage___block_26_s_y;
_q___pip_5160_1_61___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___stage___block_26_s_y : _d___pip_5160_1_61___stage___block_26_s_y;
_q___pip_5160_1_62___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___stage___block_26_s_y : _d___pip_5160_1_62___stage___block_26_s_y;
_q___pip_5160_1_63___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___stage___block_26_s_y : _d___pip_5160_1_63___stage___block_26_s_y;
_q___pip_5160_1_64___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___stage___block_26_s_y : _d___pip_5160_1_64___stage___block_26_s_y;
_q___pip_5160_1_65___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___stage___block_26_s_y : _d___pip_5160_1_65___stage___block_26_s_y;
_q___pip_5160_1_66___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___stage___block_26_s_y : _d___pip_5160_1_66___stage___block_26_s_y;
_q___pip_5160_1_67___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___stage___block_26_s_y : _d___pip_5160_1_67___stage___block_26_s_y;
_q___pip_5160_1_68___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___stage___block_26_s_y : _d___pip_5160_1_68___stage___block_26_s_y;
_q___pip_5160_1_69___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___stage___block_26_s_y : _d___pip_5160_1_69___stage___block_26_s_y;
_q___pip_5160_1_70___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___stage___block_26_s_y : _d___pip_5160_1_70___stage___block_26_s_y;
_q___pip_5160_1_71___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___stage___block_26_s_y : _d___pip_5160_1_71___stage___block_26_s_y;
_q___pip_5160_1_72___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___stage___block_26_s_y : _d___pip_5160_1_72___stage___block_26_s_y;
_q___pip_5160_1_73___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___stage___block_26_s_y : _d___pip_5160_1_73___stage___block_26_s_y;
_q___pip_5160_1_74___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___stage___block_26_s_y : _d___pip_5160_1_74___stage___block_26_s_y;
_q___pip_5160_1_75___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___stage___block_26_s_y : _d___pip_5160_1_75___stage___block_26_s_y;
_q___pip_5160_1_76___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___stage___block_26_s_y : _d___pip_5160_1_76___stage___block_26_s_y;
_q___pip_5160_1_77___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___stage___block_26_s_y : _d___pip_5160_1_77___stage___block_26_s_y;
_q___pip_5160_1_78___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___stage___block_26_s_y : _d___pip_5160_1_78___stage___block_26_s_y;
_q___pip_5160_1_79___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___stage___block_26_s_y : _d___pip_5160_1_79___stage___block_26_s_y;
_q___pip_5160_1_80___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___stage___block_26_s_y : _d___pip_5160_1_80___stage___block_26_s_y;
_q___pip_5160_1_81___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___stage___block_26_s_y : _d___pip_5160_1_81___stage___block_26_s_y;
_q___pip_5160_1_82___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___stage___block_26_s_y : _d___pip_5160_1_82___stage___block_26_s_y;
_q___pip_5160_1_83___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___stage___block_26_s_y : _d___pip_5160_1_83___stage___block_26_s_y;
_q___pip_5160_1_84___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___stage___block_26_s_y : _d___pip_5160_1_84___stage___block_26_s_y;
_q___pip_5160_1_85___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___stage___block_26_s_y : _d___pip_5160_1_85___stage___block_26_s_y;
_q___pip_5160_1_86___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___stage___block_26_s_y : _d___pip_5160_1_86___stage___block_26_s_y;
_q___pip_5160_1_87___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___stage___block_26_s_y : _d___pip_5160_1_87___stage___block_26_s_y;
_q___pip_5160_1_88___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___stage___block_26_s_y : _d___pip_5160_1_88___stage___block_26_s_y;
_q___pip_5160_1_89___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___stage___block_26_s_y : _d___pip_5160_1_89___stage___block_26_s_y;
_q___pip_5160_1_90___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___stage___block_26_s_y : _d___pip_5160_1_90___stage___block_26_s_y;
_q___pip_5160_1_91___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___stage___block_26_s_y : _d___pip_5160_1_91___stage___block_26_s_y;
_q___pip_5160_1_92___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___stage___block_26_s_y : _d___pip_5160_1_92___stage___block_26_s_y;
_q___pip_5160_1_93___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___stage___block_26_s_y : _d___pip_5160_1_93___stage___block_26_s_y;
_q___pip_5160_1_94___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___stage___block_26_s_y : _d___pip_5160_1_94___stage___block_26_s_y;
_q___pip_5160_1_95___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___stage___block_26_s_y : _d___pip_5160_1_95___stage___block_26_s_y;
_q___pip_5160_1_96___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___stage___block_26_s_y : _d___pip_5160_1_96___stage___block_26_s_y;
_q___pip_5160_1_97___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___stage___block_26_s_y : _d___pip_5160_1_97___stage___block_26_s_y;
_q___pip_5160_1_98___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___stage___block_26_s_y : _d___pip_5160_1_98___stage___block_26_s_y;
_q___pip_5160_1_99___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___stage___block_26_s_y : _d___pip_5160_1_99___stage___block_26_s_y;
_q___pip_5160_1_100___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___stage___block_26_s_y : _d___pip_5160_1_100___stage___block_26_s_y;
_q___pip_5160_1_101___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___stage___block_26_s_y : _d___pip_5160_1_101___stage___block_26_s_y;
_q___pip_5160_1_102___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___stage___block_26_s_y : _d___pip_5160_1_102___stage___block_26_s_y;
_q___pip_5160_1_103___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___stage___block_26_s_y : _d___pip_5160_1_103___stage___block_26_s_y;
_q___pip_5160_1_104___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___stage___block_26_s_y : _d___pip_5160_1_104___stage___block_26_s_y;
_q___pip_5160_1_105___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___stage___block_26_s_y : _d___pip_5160_1_105___stage___block_26_s_y;
_q___pip_5160_1_106___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___stage___block_26_s_y : _d___pip_5160_1_106___stage___block_26_s_y;
_q___pip_5160_1_107___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___stage___block_26_s_y : _d___pip_5160_1_107___stage___block_26_s_y;
_q___pip_5160_1_108___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___stage___block_26_s_y : _d___pip_5160_1_108___stage___block_26_s_y;
_q___pip_5160_1_109___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___stage___block_26_s_y : _d___pip_5160_1_109___stage___block_26_s_y;
_q___pip_5160_1_110___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___stage___block_26_s_y : _d___pip_5160_1_110___stage___block_26_s_y;
_q___pip_5160_1_111___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___stage___block_26_s_y : _d___pip_5160_1_111___stage___block_26_s_y;
_q___pip_5160_1_112___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___stage___block_26_s_y : _d___pip_5160_1_112___stage___block_26_s_y;
_q___pip_5160_1_113___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___stage___block_26_s_y : _d___pip_5160_1_113___stage___block_26_s_y;
_q___pip_5160_1_114___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___stage___block_26_s_y : _d___pip_5160_1_114___stage___block_26_s_y;
_q___pip_5160_1_115___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___stage___block_26_s_y : _d___pip_5160_1_115___stage___block_26_s_y;
_q___pip_5160_1_116___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___stage___block_26_s_y : _d___pip_5160_1_116___stage___block_26_s_y;
_q___pip_5160_1_117___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___stage___block_26_s_y : _d___pip_5160_1_117___stage___block_26_s_y;
_q___pip_5160_1_118___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___stage___block_26_s_y : _d___pip_5160_1_118___stage___block_26_s_y;
_q___pip_5160_1_119___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___stage___block_26_s_y : _d___pip_5160_1_119___stage___block_26_s_y;
_q___pip_5160_1_120___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___stage___block_26_s_y : _d___pip_5160_1_120___stage___block_26_s_y;
_q___pip_5160_1_121___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___stage___block_26_s_y : _d___pip_5160_1_121___stage___block_26_s_y;
_q___pip_5160_1_122___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___stage___block_26_s_y : _d___pip_5160_1_122___stage___block_26_s_y;
_q___pip_5160_1_123___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___stage___block_26_s_y : _d___pip_5160_1_123___stage___block_26_s_y;
_q___pip_5160_1_124___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___stage___block_26_s_y : _d___pip_5160_1_124___stage___block_26_s_y;
_q___pip_5160_1_125___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___stage___block_26_s_y : _d___pip_5160_1_125___stage___block_26_s_y;
_q___pip_5160_1_126___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___stage___block_26_s_y : _d___pip_5160_1_126___stage___block_26_s_y;
_q___pip_5160_1_127___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___stage___block_26_s_y : _d___pip_5160_1_127___stage___block_26_s_y;
_q___pip_5160_1_128___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___stage___block_26_s_y : _d___pip_5160_1_128___stage___block_26_s_y;
_q___pip_5160_1_129___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___stage___block_26_s_y : _d___pip_5160_1_129___stage___block_26_s_y;
_q___pip_5160_1_130___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___stage___block_26_s_y : _d___pip_5160_1_130___stage___block_26_s_y;
_q___pip_5160_1_131___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___stage___block_26_s_y : _d___pip_5160_1_131___stage___block_26_s_y;
_q___pip_5160_1_132___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___stage___block_26_s_y : _d___pip_5160_1_132___stage___block_26_s_y;
_q___pip_5160_1_133___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___stage___block_26_s_y : _d___pip_5160_1_133___stage___block_26_s_y;
_q___pip_5160_1_134___stage___block_26_s_y <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___stage___block_26_s_y : _d___pip_5160_1_134___stage___block_26_s_y;
_q___pip_5160_1_4___stage___block_26_s_z <= _d___pip_5160_1_4___stage___block_26_s_z;
_q___pip_5160_1_5___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_26_s_z : _d___pip_5160_1_5___stage___block_26_s_z;
_q___pip_5160_1_6___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_26_s_z : _d___pip_5160_1_6___stage___block_26_s_z;
_q___pip_5160_1_7___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___stage___block_26_s_z : _d___pip_5160_1_7___stage___block_26_s_z;
_q___pip_5160_1_8___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___stage___block_26_s_z : _d___pip_5160_1_8___stage___block_26_s_z;
_q___pip_5160_1_9___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___stage___block_26_s_z : _d___pip_5160_1_9___stage___block_26_s_z;
_q___pip_5160_1_10___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___stage___block_26_s_z : _d___pip_5160_1_10___stage___block_26_s_z;
_q___pip_5160_1_11___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___stage___block_26_s_z : _d___pip_5160_1_11___stage___block_26_s_z;
_q___pip_5160_1_12___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___stage___block_26_s_z : _d___pip_5160_1_12___stage___block_26_s_z;
_q___pip_5160_1_13___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___stage___block_26_s_z : _d___pip_5160_1_13___stage___block_26_s_z;
_q___pip_5160_1_14___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___stage___block_26_s_z : _d___pip_5160_1_14___stage___block_26_s_z;
_q___pip_5160_1_15___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___stage___block_26_s_z : _d___pip_5160_1_15___stage___block_26_s_z;
_q___pip_5160_1_16___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___stage___block_26_s_z : _d___pip_5160_1_16___stage___block_26_s_z;
_q___pip_5160_1_17___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___stage___block_26_s_z : _d___pip_5160_1_17___stage___block_26_s_z;
_q___pip_5160_1_18___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___stage___block_26_s_z : _d___pip_5160_1_18___stage___block_26_s_z;
_q___pip_5160_1_19___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___stage___block_26_s_z : _d___pip_5160_1_19___stage___block_26_s_z;
_q___pip_5160_1_20___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___stage___block_26_s_z : _d___pip_5160_1_20___stage___block_26_s_z;
_q___pip_5160_1_21___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___stage___block_26_s_z : _d___pip_5160_1_21___stage___block_26_s_z;
_q___pip_5160_1_22___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___stage___block_26_s_z : _d___pip_5160_1_22___stage___block_26_s_z;
_q___pip_5160_1_23___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___stage___block_26_s_z : _d___pip_5160_1_23___stage___block_26_s_z;
_q___pip_5160_1_24___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___stage___block_26_s_z : _d___pip_5160_1_24___stage___block_26_s_z;
_q___pip_5160_1_25___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___stage___block_26_s_z : _d___pip_5160_1_25___stage___block_26_s_z;
_q___pip_5160_1_26___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___stage___block_26_s_z : _d___pip_5160_1_26___stage___block_26_s_z;
_q___pip_5160_1_27___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___stage___block_26_s_z : _d___pip_5160_1_27___stage___block_26_s_z;
_q___pip_5160_1_28___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___stage___block_26_s_z : _d___pip_5160_1_28___stage___block_26_s_z;
_q___pip_5160_1_29___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___stage___block_26_s_z : _d___pip_5160_1_29___stage___block_26_s_z;
_q___pip_5160_1_30___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___stage___block_26_s_z : _d___pip_5160_1_30___stage___block_26_s_z;
_q___pip_5160_1_31___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___stage___block_26_s_z : _d___pip_5160_1_31___stage___block_26_s_z;
_q___pip_5160_1_32___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___stage___block_26_s_z : _d___pip_5160_1_32___stage___block_26_s_z;
_q___pip_5160_1_33___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___stage___block_26_s_z : _d___pip_5160_1_33___stage___block_26_s_z;
_q___pip_5160_1_34___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___stage___block_26_s_z : _d___pip_5160_1_34___stage___block_26_s_z;
_q___pip_5160_1_35___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___stage___block_26_s_z : _d___pip_5160_1_35___stage___block_26_s_z;
_q___pip_5160_1_36___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___stage___block_26_s_z : _d___pip_5160_1_36___stage___block_26_s_z;
_q___pip_5160_1_37___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___stage___block_26_s_z : _d___pip_5160_1_37___stage___block_26_s_z;
_q___pip_5160_1_38___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___stage___block_26_s_z : _d___pip_5160_1_38___stage___block_26_s_z;
_q___pip_5160_1_39___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___stage___block_26_s_z : _d___pip_5160_1_39___stage___block_26_s_z;
_q___pip_5160_1_40___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___stage___block_26_s_z : _d___pip_5160_1_40___stage___block_26_s_z;
_q___pip_5160_1_41___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___stage___block_26_s_z : _d___pip_5160_1_41___stage___block_26_s_z;
_q___pip_5160_1_42___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___stage___block_26_s_z : _d___pip_5160_1_42___stage___block_26_s_z;
_q___pip_5160_1_43___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___stage___block_26_s_z : _d___pip_5160_1_43___stage___block_26_s_z;
_q___pip_5160_1_44___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___stage___block_26_s_z : _d___pip_5160_1_44___stage___block_26_s_z;
_q___pip_5160_1_45___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___stage___block_26_s_z : _d___pip_5160_1_45___stage___block_26_s_z;
_q___pip_5160_1_46___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___stage___block_26_s_z : _d___pip_5160_1_46___stage___block_26_s_z;
_q___pip_5160_1_47___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___stage___block_26_s_z : _d___pip_5160_1_47___stage___block_26_s_z;
_q___pip_5160_1_48___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___stage___block_26_s_z : _d___pip_5160_1_48___stage___block_26_s_z;
_q___pip_5160_1_49___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___stage___block_26_s_z : _d___pip_5160_1_49___stage___block_26_s_z;
_q___pip_5160_1_50___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___stage___block_26_s_z : _d___pip_5160_1_50___stage___block_26_s_z;
_q___pip_5160_1_51___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___stage___block_26_s_z : _d___pip_5160_1_51___stage___block_26_s_z;
_q___pip_5160_1_52___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___stage___block_26_s_z : _d___pip_5160_1_52___stage___block_26_s_z;
_q___pip_5160_1_53___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___stage___block_26_s_z : _d___pip_5160_1_53___stage___block_26_s_z;
_q___pip_5160_1_54___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___stage___block_26_s_z : _d___pip_5160_1_54___stage___block_26_s_z;
_q___pip_5160_1_55___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___stage___block_26_s_z : _d___pip_5160_1_55___stage___block_26_s_z;
_q___pip_5160_1_56___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___stage___block_26_s_z : _d___pip_5160_1_56___stage___block_26_s_z;
_q___pip_5160_1_57___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___stage___block_26_s_z : _d___pip_5160_1_57___stage___block_26_s_z;
_q___pip_5160_1_58___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___stage___block_26_s_z : _d___pip_5160_1_58___stage___block_26_s_z;
_q___pip_5160_1_59___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___stage___block_26_s_z : _d___pip_5160_1_59___stage___block_26_s_z;
_q___pip_5160_1_60___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___stage___block_26_s_z : _d___pip_5160_1_60___stage___block_26_s_z;
_q___pip_5160_1_61___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___stage___block_26_s_z : _d___pip_5160_1_61___stage___block_26_s_z;
_q___pip_5160_1_62___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___stage___block_26_s_z : _d___pip_5160_1_62___stage___block_26_s_z;
_q___pip_5160_1_63___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___stage___block_26_s_z : _d___pip_5160_1_63___stage___block_26_s_z;
_q___pip_5160_1_64___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___stage___block_26_s_z : _d___pip_5160_1_64___stage___block_26_s_z;
_q___pip_5160_1_65___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___stage___block_26_s_z : _d___pip_5160_1_65___stage___block_26_s_z;
_q___pip_5160_1_66___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___stage___block_26_s_z : _d___pip_5160_1_66___stage___block_26_s_z;
_q___pip_5160_1_67___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___stage___block_26_s_z : _d___pip_5160_1_67___stage___block_26_s_z;
_q___pip_5160_1_68___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___stage___block_26_s_z : _d___pip_5160_1_68___stage___block_26_s_z;
_q___pip_5160_1_69___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___stage___block_26_s_z : _d___pip_5160_1_69___stage___block_26_s_z;
_q___pip_5160_1_70___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___stage___block_26_s_z : _d___pip_5160_1_70___stage___block_26_s_z;
_q___pip_5160_1_71___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___stage___block_26_s_z : _d___pip_5160_1_71___stage___block_26_s_z;
_q___pip_5160_1_72___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___stage___block_26_s_z : _d___pip_5160_1_72___stage___block_26_s_z;
_q___pip_5160_1_73___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___stage___block_26_s_z : _d___pip_5160_1_73___stage___block_26_s_z;
_q___pip_5160_1_74___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___stage___block_26_s_z : _d___pip_5160_1_74___stage___block_26_s_z;
_q___pip_5160_1_75___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___stage___block_26_s_z : _d___pip_5160_1_75___stage___block_26_s_z;
_q___pip_5160_1_76___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___stage___block_26_s_z : _d___pip_5160_1_76___stage___block_26_s_z;
_q___pip_5160_1_77___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___stage___block_26_s_z : _d___pip_5160_1_77___stage___block_26_s_z;
_q___pip_5160_1_78___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___stage___block_26_s_z : _d___pip_5160_1_78___stage___block_26_s_z;
_q___pip_5160_1_79___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___stage___block_26_s_z : _d___pip_5160_1_79___stage___block_26_s_z;
_q___pip_5160_1_80___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___stage___block_26_s_z : _d___pip_5160_1_80___stage___block_26_s_z;
_q___pip_5160_1_81___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___stage___block_26_s_z : _d___pip_5160_1_81___stage___block_26_s_z;
_q___pip_5160_1_82___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___stage___block_26_s_z : _d___pip_5160_1_82___stage___block_26_s_z;
_q___pip_5160_1_83___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___stage___block_26_s_z : _d___pip_5160_1_83___stage___block_26_s_z;
_q___pip_5160_1_84___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___stage___block_26_s_z : _d___pip_5160_1_84___stage___block_26_s_z;
_q___pip_5160_1_85___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___stage___block_26_s_z : _d___pip_5160_1_85___stage___block_26_s_z;
_q___pip_5160_1_86___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___stage___block_26_s_z : _d___pip_5160_1_86___stage___block_26_s_z;
_q___pip_5160_1_87___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___stage___block_26_s_z : _d___pip_5160_1_87___stage___block_26_s_z;
_q___pip_5160_1_88___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___stage___block_26_s_z : _d___pip_5160_1_88___stage___block_26_s_z;
_q___pip_5160_1_89___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___stage___block_26_s_z : _d___pip_5160_1_89___stage___block_26_s_z;
_q___pip_5160_1_90___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___stage___block_26_s_z : _d___pip_5160_1_90___stage___block_26_s_z;
_q___pip_5160_1_91___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___stage___block_26_s_z : _d___pip_5160_1_91___stage___block_26_s_z;
_q___pip_5160_1_92___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___stage___block_26_s_z : _d___pip_5160_1_92___stage___block_26_s_z;
_q___pip_5160_1_93___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___stage___block_26_s_z : _d___pip_5160_1_93___stage___block_26_s_z;
_q___pip_5160_1_94___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___stage___block_26_s_z : _d___pip_5160_1_94___stage___block_26_s_z;
_q___pip_5160_1_95___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___stage___block_26_s_z : _d___pip_5160_1_95___stage___block_26_s_z;
_q___pip_5160_1_96___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___stage___block_26_s_z : _d___pip_5160_1_96___stage___block_26_s_z;
_q___pip_5160_1_97___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___stage___block_26_s_z : _d___pip_5160_1_97___stage___block_26_s_z;
_q___pip_5160_1_98___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___stage___block_26_s_z : _d___pip_5160_1_98___stage___block_26_s_z;
_q___pip_5160_1_99___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___stage___block_26_s_z : _d___pip_5160_1_99___stage___block_26_s_z;
_q___pip_5160_1_100___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___stage___block_26_s_z : _d___pip_5160_1_100___stage___block_26_s_z;
_q___pip_5160_1_101___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___stage___block_26_s_z : _d___pip_5160_1_101___stage___block_26_s_z;
_q___pip_5160_1_102___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___stage___block_26_s_z : _d___pip_5160_1_102___stage___block_26_s_z;
_q___pip_5160_1_103___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___stage___block_26_s_z : _d___pip_5160_1_103___stage___block_26_s_z;
_q___pip_5160_1_104___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___stage___block_26_s_z : _d___pip_5160_1_104___stage___block_26_s_z;
_q___pip_5160_1_105___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___stage___block_26_s_z : _d___pip_5160_1_105___stage___block_26_s_z;
_q___pip_5160_1_106___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___stage___block_26_s_z : _d___pip_5160_1_106___stage___block_26_s_z;
_q___pip_5160_1_107___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___stage___block_26_s_z : _d___pip_5160_1_107___stage___block_26_s_z;
_q___pip_5160_1_108___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___stage___block_26_s_z : _d___pip_5160_1_108___stage___block_26_s_z;
_q___pip_5160_1_109___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___stage___block_26_s_z : _d___pip_5160_1_109___stage___block_26_s_z;
_q___pip_5160_1_110___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___stage___block_26_s_z : _d___pip_5160_1_110___stage___block_26_s_z;
_q___pip_5160_1_111___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___stage___block_26_s_z : _d___pip_5160_1_111___stage___block_26_s_z;
_q___pip_5160_1_112___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___stage___block_26_s_z : _d___pip_5160_1_112___stage___block_26_s_z;
_q___pip_5160_1_113___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___stage___block_26_s_z : _d___pip_5160_1_113___stage___block_26_s_z;
_q___pip_5160_1_114___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___stage___block_26_s_z : _d___pip_5160_1_114___stage___block_26_s_z;
_q___pip_5160_1_115___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___stage___block_26_s_z : _d___pip_5160_1_115___stage___block_26_s_z;
_q___pip_5160_1_116___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___stage___block_26_s_z : _d___pip_5160_1_116___stage___block_26_s_z;
_q___pip_5160_1_117___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___stage___block_26_s_z : _d___pip_5160_1_117___stage___block_26_s_z;
_q___pip_5160_1_118___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___stage___block_26_s_z : _d___pip_5160_1_118___stage___block_26_s_z;
_q___pip_5160_1_119___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___stage___block_26_s_z : _d___pip_5160_1_119___stage___block_26_s_z;
_q___pip_5160_1_120___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___stage___block_26_s_z : _d___pip_5160_1_120___stage___block_26_s_z;
_q___pip_5160_1_121___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___stage___block_26_s_z : _d___pip_5160_1_121___stage___block_26_s_z;
_q___pip_5160_1_122___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___stage___block_26_s_z : _d___pip_5160_1_122___stage___block_26_s_z;
_q___pip_5160_1_123___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___stage___block_26_s_z : _d___pip_5160_1_123___stage___block_26_s_z;
_q___pip_5160_1_124___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___stage___block_26_s_z : _d___pip_5160_1_124___stage___block_26_s_z;
_q___pip_5160_1_125___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___stage___block_26_s_z : _d___pip_5160_1_125___stage___block_26_s_z;
_q___pip_5160_1_126___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___stage___block_26_s_z : _d___pip_5160_1_126___stage___block_26_s_z;
_q___pip_5160_1_127___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___stage___block_26_s_z : _d___pip_5160_1_127___stage___block_26_s_z;
_q___pip_5160_1_128___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___stage___block_26_s_z : _d___pip_5160_1_128___stage___block_26_s_z;
_q___pip_5160_1_129___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___stage___block_26_s_z : _d___pip_5160_1_129___stage___block_26_s_z;
_q___pip_5160_1_130___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___stage___block_26_s_z : _d___pip_5160_1_130___stage___block_26_s_z;
_q___pip_5160_1_131___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___stage___block_26_s_z : _d___pip_5160_1_131___stage___block_26_s_z;
_q___pip_5160_1_132___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___stage___block_26_s_z : _d___pip_5160_1_132___stage___block_26_s_z;
_q___pip_5160_1_133___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___stage___block_26_s_z : _d___pip_5160_1_133___stage___block_26_s_z;
_q___pip_5160_1_134___stage___block_26_s_z <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___stage___block_26_s_z : _d___pip_5160_1_134___stage___block_26_s_z;
_q___pip_5160_1_4___stage___block_26_v_x <= _d___pip_5160_1_4___stage___block_26_v_x;
_q___pip_5160_1_5___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_26_v_x : _d___pip_5160_1_5___stage___block_26_v_x;
_q___pip_5160_1_6___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_26_v_x : _d___pip_5160_1_6___stage___block_26_v_x;
_q___pip_5160_1_7___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___stage___block_26_v_x : _d___pip_5160_1_7___stage___block_26_v_x;
_q___pip_5160_1_8___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___stage___block_26_v_x : _d___pip_5160_1_8___stage___block_26_v_x;
_q___pip_5160_1_9___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___stage___block_26_v_x : _d___pip_5160_1_9___stage___block_26_v_x;
_q___pip_5160_1_10___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___stage___block_26_v_x : _d___pip_5160_1_10___stage___block_26_v_x;
_q___pip_5160_1_11___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___stage___block_26_v_x : _d___pip_5160_1_11___stage___block_26_v_x;
_q___pip_5160_1_12___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___stage___block_26_v_x : _d___pip_5160_1_12___stage___block_26_v_x;
_q___pip_5160_1_13___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___stage___block_26_v_x : _d___pip_5160_1_13___stage___block_26_v_x;
_q___pip_5160_1_14___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___stage___block_26_v_x : _d___pip_5160_1_14___stage___block_26_v_x;
_q___pip_5160_1_15___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___stage___block_26_v_x : _d___pip_5160_1_15___stage___block_26_v_x;
_q___pip_5160_1_16___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___stage___block_26_v_x : _d___pip_5160_1_16___stage___block_26_v_x;
_q___pip_5160_1_17___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___stage___block_26_v_x : _d___pip_5160_1_17___stage___block_26_v_x;
_q___pip_5160_1_18___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___stage___block_26_v_x : _d___pip_5160_1_18___stage___block_26_v_x;
_q___pip_5160_1_19___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___stage___block_26_v_x : _d___pip_5160_1_19___stage___block_26_v_x;
_q___pip_5160_1_20___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___stage___block_26_v_x : _d___pip_5160_1_20___stage___block_26_v_x;
_q___pip_5160_1_21___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___stage___block_26_v_x : _d___pip_5160_1_21___stage___block_26_v_x;
_q___pip_5160_1_22___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___stage___block_26_v_x : _d___pip_5160_1_22___stage___block_26_v_x;
_q___pip_5160_1_23___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___stage___block_26_v_x : _d___pip_5160_1_23___stage___block_26_v_x;
_q___pip_5160_1_24___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___stage___block_26_v_x : _d___pip_5160_1_24___stage___block_26_v_x;
_q___pip_5160_1_25___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___stage___block_26_v_x : _d___pip_5160_1_25___stage___block_26_v_x;
_q___pip_5160_1_26___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___stage___block_26_v_x : _d___pip_5160_1_26___stage___block_26_v_x;
_q___pip_5160_1_27___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___stage___block_26_v_x : _d___pip_5160_1_27___stage___block_26_v_x;
_q___pip_5160_1_28___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___stage___block_26_v_x : _d___pip_5160_1_28___stage___block_26_v_x;
_q___pip_5160_1_29___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___stage___block_26_v_x : _d___pip_5160_1_29___stage___block_26_v_x;
_q___pip_5160_1_30___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___stage___block_26_v_x : _d___pip_5160_1_30___stage___block_26_v_x;
_q___pip_5160_1_31___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___stage___block_26_v_x : _d___pip_5160_1_31___stage___block_26_v_x;
_q___pip_5160_1_32___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___stage___block_26_v_x : _d___pip_5160_1_32___stage___block_26_v_x;
_q___pip_5160_1_33___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___stage___block_26_v_x : _d___pip_5160_1_33___stage___block_26_v_x;
_q___pip_5160_1_34___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___stage___block_26_v_x : _d___pip_5160_1_34___stage___block_26_v_x;
_q___pip_5160_1_35___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___stage___block_26_v_x : _d___pip_5160_1_35___stage___block_26_v_x;
_q___pip_5160_1_36___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___stage___block_26_v_x : _d___pip_5160_1_36___stage___block_26_v_x;
_q___pip_5160_1_37___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___stage___block_26_v_x : _d___pip_5160_1_37___stage___block_26_v_x;
_q___pip_5160_1_38___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___stage___block_26_v_x : _d___pip_5160_1_38___stage___block_26_v_x;
_q___pip_5160_1_39___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___stage___block_26_v_x : _d___pip_5160_1_39___stage___block_26_v_x;
_q___pip_5160_1_40___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___stage___block_26_v_x : _d___pip_5160_1_40___stage___block_26_v_x;
_q___pip_5160_1_41___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___stage___block_26_v_x : _d___pip_5160_1_41___stage___block_26_v_x;
_q___pip_5160_1_42___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___stage___block_26_v_x : _d___pip_5160_1_42___stage___block_26_v_x;
_q___pip_5160_1_43___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___stage___block_26_v_x : _d___pip_5160_1_43___stage___block_26_v_x;
_q___pip_5160_1_44___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___stage___block_26_v_x : _d___pip_5160_1_44___stage___block_26_v_x;
_q___pip_5160_1_45___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___stage___block_26_v_x : _d___pip_5160_1_45___stage___block_26_v_x;
_q___pip_5160_1_46___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___stage___block_26_v_x : _d___pip_5160_1_46___stage___block_26_v_x;
_q___pip_5160_1_47___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___stage___block_26_v_x : _d___pip_5160_1_47___stage___block_26_v_x;
_q___pip_5160_1_48___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___stage___block_26_v_x : _d___pip_5160_1_48___stage___block_26_v_x;
_q___pip_5160_1_49___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___stage___block_26_v_x : _d___pip_5160_1_49___stage___block_26_v_x;
_q___pip_5160_1_50___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___stage___block_26_v_x : _d___pip_5160_1_50___stage___block_26_v_x;
_q___pip_5160_1_51___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___stage___block_26_v_x : _d___pip_5160_1_51___stage___block_26_v_x;
_q___pip_5160_1_52___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___stage___block_26_v_x : _d___pip_5160_1_52___stage___block_26_v_x;
_q___pip_5160_1_53___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___stage___block_26_v_x : _d___pip_5160_1_53___stage___block_26_v_x;
_q___pip_5160_1_54___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___stage___block_26_v_x : _d___pip_5160_1_54___stage___block_26_v_x;
_q___pip_5160_1_55___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___stage___block_26_v_x : _d___pip_5160_1_55___stage___block_26_v_x;
_q___pip_5160_1_56___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___stage___block_26_v_x : _d___pip_5160_1_56___stage___block_26_v_x;
_q___pip_5160_1_57___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___stage___block_26_v_x : _d___pip_5160_1_57___stage___block_26_v_x;
_q___pip_5160_1_58___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___stage___block_26_v_x : _d___pip_5160_1_58___stage___block_26_v_x;
_q___pip_5160_1_59___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___stage___block_26_v_x : _d___pip_5160_1_59___stage___block_26_v_x;
_q___pip_5160_1_60___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___stage___block_26_v_x : _d___pip_5160_1_60___stage___block_26_v_x;
_q___pip_5160_1_61___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___stage___block_26_v_x : _d___pip_5160_1_61___stage___block_26_v_x;
_q___pip_5160_1_62___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___stage___block_26_v_x : _d___pip_5160_1_62___stage___block_26_v_x;
_q___pip_5160_1_63___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___stage___block_26_v_x : _d___pip_5160_1_63___stage___block_26_v_x;
_q___pip_5160_1_64___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___stage___block_26_v_x : _d___pip_5160_1_64___stage___block_26_v_x;
_q___pip_5160_1_65___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___stage___block_26_v_x : _d___pip_5160_1_65___stage___block_26_v_x;
_q___pip_5160_1_66___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___stage___block_26_v_x : _d___pip_5160_1_66___stage___block_26_v_x;
_q___pip_5160_1_67___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___stage___block_26_v_x : _d___pip_5160_1_67___stage___block_26_v_x;
_q___pip_5160_1_68___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___stage___block_26_v_x : _d___pip_5160_1_68___stage___block_26_v_x;
_q___pip_5160_1_69___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___stage___block_26_v_x : _d___pip_5160_1_69___stage___block_26_v_x;
_q___pip_5160_1_70___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___stage___block_26_v_x : _d___pip_5160_1_70___stage___block_26_v_x;
_q___pip_5160_1_71___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___stage___block_26_v_x : _d___pip_5160_1_71___stage___block_26_v_x;
_q___pip_5160_1_72___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___stage___block_26_v_x : _d___pip_5160_1_72___stage___block_26_v_x;
_q___pip_5160_1_73___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___stage___block_26_v_x : _d___pip_5160_1_73___stage___block_26_v_x;
_q___pip_5160_1_74___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___stage___block_26_v_x : _d___pip_5160_1_74___stage___block_26_v_x;
_q___pip_5160_1_75___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___stage___block_26_v_x : _d___pip_5160_1_75___stage___block_26_v_x;
_q___pip_5160_1_76___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___stage___block_26_v_x : _d___pip_5160_1_76___stage___block_26_v_x;
_q___pip_5160_1_77___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___stage___block_26_v_x : _d___pip_5160_1_77___stage___block_26_v_x;
_q___pip_5160_1_78___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___stage___block_26_v_x : _d___pip_5160_1_78___stage___block_26_v_x;
_q___pip_5160_1_79___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___stage___block_26_v_x : _d___pip_5160_1_79___stage___block_26_v_x;
_q___pip_5160_1_80___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___stage___block_26_v_x : _d___pip_5160_1_80___stage___block_26_v_x;
_q___pip_5160_1_81___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___stage___block_26_v_x : _d___pip_5160_1_81___stage___block_26_v_x;
_q___pip_5160_1_82___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___stage___block_26_v_x : _d___pip_5160_1_82___stage___block_26_v_x;
_q___pip_5160_1_83___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___stage___block_26_v_x : _d___pip_5160_1_83___stage___block_26_v_x;
_q___pip_5160_1_84___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___stage___block_26_v_x : _d___pip_5160_1_84___stage___block_26_v_x;
_q___pip_5160_1_85___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___stage___block_26_v_x : _d___pip_5160_1_85___stage___block_26_v_x;
_q___pip_5160_1_86___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___stage___block_26_v_x : _d___pip_5160_1_86___stage___block_26_v_x;
_q___pip_5160_1_87___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___stage___block_26_v_x : _d___pip_5160_1_87___stage___block_26_v_x;
_q___pip_5160_1_88___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___stage___block_26_v_x : _d___pip_5160_1_88___stage___block_26_v_x;
_q___pip_5160_1_89___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___stage___block_26_v_x : _d___pip_5160_1_89___stage___block_26_v_x;
_q___pip_5160_1_90___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___stage___block_26_v_x : _d___pip_5160_1_90___stage___block_26_v_x;
_q___pip_5160_1_91___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___stage___block_26_v_x : _d___pip_5160_1_91___stage___block_26_v_x;
_q___pip_5160_1_92___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___stage___block_26_v_x : _d___pip_5160_1_92___stage___block_26_v_x;
_q___pip_5160_1_93___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___stage___block_26_v_x : _d___pip_5160_1_93___stage___block_26_v_x;
_q___pip_5160_1_94___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___stage___block_26_v_x : _d___pip_5160_1_94___stage___block_26_v_x;
_q___pip_5160_1_95___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___stage___block_26_v_x : _d___pip_5160_1_95___stage___block_26_v_x;
_q___pip_5160_1_96___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___stage___block_26_v_x : _d___pip_5160_1_96___stage___block_26_v_x;
_q___pip_5160_1_97___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___stage___block_26_v_x : _d___pip_5160_1_97___stage___block_26_v_x;
_q___pip_5160_1_98___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___stage___block_26_v_x : _d___pip_5160_1_98___stage___block_26_v_x;
_q___pip_5160_1_99___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___stage___block_26_v_x : _d___pip_5160_1_99___stage___block_26_v_x;
_q___pip_5160_1_100___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___stage___block_26_v_x : _d___pip_5160_1_100___stage___block_26_v_x;
_q___pip_5160_1_101___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___stage___block_26_v_x : _d___pip_5160_1_101___stage___block_26_v_x;
_q___pip_5160_1_102___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___stage___block_26_v_x : _d___pip_5160_1_102___stage___block_26_v_x;
_q___pip_5160_1_103___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___stage___block_26_v_x : _d___pip_5160_1_103___stage___block_26_v_x;
_q___pip_5160_1_104___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___stage___block_26_v_x : _d___pip_5160_1_104___stage___block_26_v_x;
_q___pip_5160_1_105___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___stage___block_26_v_x : _d___pip_5160_1_105___stage___block_26_v_x;
_q___pip_5160_1_106___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___stage___block_26_v_x : _d___pip_5160_1_106___stage___block_26_v_x;
_q___pip_5160_1_107___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___stage___block_26_v_x : _d___pip_5160_1_107___stage___block_26_v_x;
_q___pip_5160_1_108___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___stage___block_26_v_x : _d___pip_5160_1_108___stage___block_26_v_x;
_q___pip_5160_1_109___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___stage___block_26_v_x : _d___pip_5160_1_109___stage___block_26_v_x;
_q___pip_5160_1_110___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___stage___block_26_v_x : _d___pip_5160_1_110___stage___block_26_v_x;
_q___pip_5160_1_111___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___stage___block_26_v_x : _d___pip_5160_1_111___stage___block_26_v_x;
_q___pip_5160_1_112___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___stage___block_26_v_x : _d___pip_5160_1_112___stage___block_26_v_x;
_q___pip_5160_1_113___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___stage___block_26_v_x : _d___pip_5160_1_113___stage___block_26_v_x;
_q___pip_5160_1_114___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___stage___block_26_v_x : _d___pip_5160_1_114___stage___block_26_v_x;
_q___pip_5160_1_115___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___stage___block_26_v_x : _d___pip_5160_1_115___stage___block_26_v_x;
_q___pip_5160_1_116___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___stage___block_26_v_x : _d___pip_5160_1_116___stage___block_26_v_x;
_q___pip_5160_1_117___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___stage___block_26_v_x : _d___pip_5160_1_117___stage___block_26_v_x;
_q___pip_5160_1_118___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___stage___block_26_v_x : _d___pip_5160_1_118___stage___block_26_v_x;
_q___pip_5160_1_119___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___stage___block_26_v_x : _d___pip_5160_1_119___stage___block_26_v_x;
_q___pip_5160_1_120___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___stage___block_26_v_x : _d___pip_5160_1_120___stage___block_26_v_x;
_q___pip_5160_1_121___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___stage___block_26_v_x : _d___pip_5160_1_121___stage___block_26_v_x;
_q___pip_5160_1_122___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___stage___block_26_v_x : _d___pip_5160_1_122___stage___block_26_v_x;
_q___pip_5160_1_123___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___stage___block_26_v_x : _d___pip_5160_1_123___stage___block_26_v_x;
_q___pip_5160_1_124___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___stage___block_26_v_x : _d___pip_5160_1_124___stage___block_26_v_x;
_q___pip_5160_1_125___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___stage___block_26_v_x : _d___pip_5160_1_125___stage___block_26_v_x;
_q___pip_5160_1_126___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___stage___block_26_v_x : _d___pip_5160_1_126___stage___block_26_v_x;
_q___pip_5160_1_127___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___stage___block_26_v_x : _d___pip_5160_1_127___stage___block_26_v_x;
_q___pip_5160_1_128___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___stage___block_26_v_x : _d___pip_5160_1_128___stage___block_26_v_x;
_q___pip_5160_1_129___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___stage___block_26_v_x : _d___pip_5160_1_129___stage___block_26_v_x;
_q___pip_5160_1_130___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___stage___block_26_v_x : _d___pip_5160_1_130___stage___block_26_v_x;
_q___pip_5160_1_131___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___stage___block_26_v_x : _d___pip_5160_1_131___stage___block_26_v_x;
_q___pip_5160_1_132___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___stage___block_26_v_x : _d___pip_5160_1_132___stage___block_26_v_x;
_q___pip_5160_1_133___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___stage___block_26_v_x : _d___pip_5160_1_133___stage___block_26_v_x;
_q___pip_5160_1_134___stage___block_26_v_x <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___stage___block_26_v_x : _d___pip_5160_1_134___stage___block_26_v_x;
_q___pip_5160_1_4___stage___block_26_v_y <= _d___pip_5160_1_4___stage___block_26_v_y;
_q___pip_5160_1_5___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_26_v_y : _d___pip_5160_1_5___stage___block_26_v_y;
_q___pip_5160_1_6___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_26_v_y : _d___pip_5160_1_6___stage___block_26_v_y;
_q___pip_5160_1_7___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___stage___block_26_v_y : _d___pip_5160_1_7___stage___block_26_v_y;
_q___pip_5160_1_8___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___stage___block_26_v_y : _d___pip_5160_1_8___stage___block_26_v_y;
_q___pip_5160_1_9___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___stage___block_26_v_y : _d___pip_5160_1_9___stage___block_26_v_y;
_q___pip_5160_1_10___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___stage___block_26_v_y : _d___pip_5160_1_10___stage___block_26_v_y;
_q___pip_5160_1_11___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___stage___block_26_v_y : _d___pip_5160_1_11___stage___block_26_v_y;
_q___pip_5160_1_12___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___stage___block_26_v_y : _d___pip_5160_1_12___stage___block_26_v_y;
_q___pip_5160_1_13___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___stage___block_26_v_y : _d___pip_5160_1_13___stage___block_26_v_y;
_q___pip_5160_1_14___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___stage___block_26_v_y : _d___pip_5160_1_14___stage___block_26_v_y;
_q___pip_5160_1_15___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___stage___block_26_v_y : _d___pip_5160_1_15___stage___block_26_v_y;
_q___pip_5160_1_16___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___stage___block_26_v_y : _d___pip_5160_1_16___stage___block_26_v_y;
_q___pip_5160_1_17___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___stage___block_26_v_y : _d___pip_5160_1_17___stage___block_26_v_y;
_q___pip_5160_1_18___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___stage___block_26_v_y : _d___pip_5160_1_18___stage___block_26_v_y;
_q___pip_5160_1_19___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___stage___block_26_v_y : _d___pip_5160_1_19___stage___block_26_v_y;
_q___pip_5160_1_20___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___stage___block_26_v_y : _d___pip_5160_1_20___stage___block_26_v_y;
_q___pip_5160_1_21___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___stage___block_26_v_y : _d___pip_5160_1_21___stage___block_26_v_y;
_q___pip_5160_1_22___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___stage___block_26_v_y : _d___pip_5160_1_22___stage___block_26_v_y;
_q___pip_5160_1_23___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___stage___block_26_v_y : _d___pip_5160_1_23___stage___block_26_v_y;
_q___pip_5160_1_24___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___stage___block_26_v_y : _d___pip_5160_1_24___stage___block_26_v_y;
_q___pip_5160_1_25___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___stage___block_26_v_y : _d___pip_5160_1_25___stage___block_26_v_y;
_q___pip_5160_1_26___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___stage___block_26_v_y : _d___pip_5160_1_26___stage___block_26_v_y;
_q___pip_5160_1_27___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___stage___block_26_v_y : _d___pip_5160_1_27___stage___block_26_v_y;
_q___pip_5160_1_28___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___stage___block_26_v_y : _d___pip_5160_1_28___stage___block_26_v_y;
_q___pip_5160_1_29___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___stage___block_26_v_y : _d___pip_5160_1_29___stage___block_26_v_y;
_q___pip_5160_1_30___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___stage___block_26_v_y : _d___pip_5160_1_30___stage___block_26_v_y;
_q___pip_5160_1_31___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___stage___block_26_v_y : _d___pip_5160_1_31___stage___block_26_v_y;
_q___pip_5160_1_32___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___stage___block_26_v_y : _d___pip_5160_1_32___stage___block_26_v_y;
_q___pip_5160_1_33___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___stage___block_26_v_y : _d___pip_5160_1_33___stage___block_26_v_y;
_q___pip_5160_1_34___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___stage___block_26_v_y : _d___pip_5160_1_34___stage___block_26_v_y;
_q___pip_5160_1_35___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___stage___block_26_v_y : _d___pip_5160_1_35___stage___block_26_v_y;
_q___pip_5160_1_36___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___stage___block_26_v_y : _d___pip_5160_1_36___stage___block_26_v_y;
_q___pip_5160_1_37___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___stage___block_26_v_y : _d___pip_5160_1_37___stage___block_26_v_y;
_q___pip_5160_1_38___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___stage___block_26_v_y : _d___pip_5160_1_38___stage___block_26_v_y;
_q___pip_5160_1_39___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___stage___block_26_v_y : _d___pip_5160_1_39___stage___block_26_v_y;
_q___pip_5160_1_40___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___stage___block_26_v_y : _d___pip_5160_1_40___stage___block_26_v_y;
_q___pip_5160_1_41___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___stage___block_26_v_y : _d___pip_5160_1_41___stage___block_26_v_y;
_q___pip_5160_1_42___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___stage___block_26_v_y : _d___pip_5160_1_42___stage___block_26_v_y;
_q___pip_5160_1_43___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___stage___block_26_v_y : _d___pip_5160_1_43___stage___block_26_v_y;
_q___pip_5160_1_44___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___stage___block_26_v_y : _d___pip_5160_1_44___stage___block_26_v_y;
_q___pip_5160_1_45___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___stage___block_26_v_y : _d___pip_5160_1_45___stage___block_26_v_y;
_q___pip_5160_1_46___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___stage___block_26_v_y : _d___pip_5160_1_46___stage___block_26_v_y;
_q___pip_5160_1_47___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___stage___block_26_v_y : _d___pip_5160_1_47___stage___block_26_v_y;
_q___pip_5160_1_48___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___stage___block_26_v_y : _d___pip_5160_1_48___stage___block_26_v_y;
_q___pip_5160_1_49___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___stage___block_26_v_y : _d___pip_5160_1_49___stage___block_26_v_y;
_q___pip_5160_1_50___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___stage___block_26_v_y : _d___pip_5160_1_50___stage___block_26_v_y;
_q___pip_5160_1_51___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___stage___block_26_v_y : _d___pip_5160_1_51___stage___block_26_v_y;
_q___pip_5160_1_52___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___stage___block_26_v_y : _d___pip_5160_1_52___stage___block_26_v_y;
_q___pip_5160_1_53___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___stage___block_26_v_y : _d___pip_5160_1_53___stage___block_26_v_y;
_q___pip_5160_1_54___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___stage___block_26_v_y : _d___pip_5160_1_54___stage___block_26_v_y;
_q___pip_5160_1_55___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___stage___block_26_v_y : _d___pip_5160_1_55___stage___block_26_v_y;
_q___pip_5160_1_56___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___stage___block_26_v_y : _d___pip_5160_1_56___stage___block_26_v_y;
_q___pip_5160_1_57___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___stage___block_26_v_y : _d___pip_5160_1_57___stage___block_26_v_y;
_q___pip_5160_1_58___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___stage___block_26_v_y : _d___pip_5160_1_58___stage___block_26_v_y;
_q___pip_5160_1_59___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___stage___block_26_v_y : _d___pip_5160_1_59___stage___block_26_v_y;
_q___pip_5160_1_60___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___stage___block_26_v_y : _d___pip_5160_1_60___stage___block_26_v_y;
_q___pip_5160_1_61___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___stage___block_26_v_y : _d___pip_5160_1_61___stage___block_26_v_y;
_q___pip_5160_1_62___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___stage___block_26_v_y : _d___pip_5160_1_62___stage___block_26_v_y;
_q___pip_5160_1_63___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___stage___block_26_v_y : _d___pip_5160_1_63___stage___block_26_v_y;
_q___pip_5160_1_64___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___stage___block_26_v_y : _d___pip_5160_1_64___stage___block_26_v_y;
_q___pip_5160_1_65___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___stage___block_26_v_y : _d___pip_5160_1_65___stage___block_26_v_y;
_q___pip_5160_1_66___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___stage___block_26_v_y : _d___pip_5160_1_66___stage___block_26_v_y;
_q___pip_5160_1_67___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___stage___block_26_v_y : _d___pip_5160_1_67___stage___block_26_v_y;
_q___pip_5160_1_68___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___stage___block_26_v_y : _d___pip_5160_1_68___stage___block_26_v_y;
_q___pip_5160_1_69___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___stage___block_26_v_y : _d___pip_5160_1_69___stage___block_26_v_y;
_q___pip_5160_1_70___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___stage___block_26_v_y : _d___pip_5160_1_70___stage___block_26_v_y;
_q___pip_5160_1_71___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___stage___block_26_v_y : _d___pip_5160_1_71___stage___block_26_v_y;
_q___pip_5160_1_72___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___stage___block_26_v_y : _d___pip_5160_1_72___stage___block_26_v_y;
_q___pip_5160_1_73___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___stage___block_26_v_y : _d___pip_5160_1_73___stage___block_26_v_y;
_q___pip_5160_1_74___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___stage___block_26_v_y : _d___pip_5160_1_74___stage___block_26_v_y;
_q___pip_5160_1_75___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___stage___block_26_v_y : _d___pip_5160_1_75___stage___block_26_v_y;
_q___pip_5160_1_76___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___stage___block_26_v_y : _d___pip_5160_1_76___stage___block_26_v_y;
_q___pip_5160_1_77___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___stage___block_26_v_y : _d___pip_5160_1_77___stage___block_26_v_y;
_q___pip_5160_1_78___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___stage___block_26_v_y : _d___pip_5160_1_78___stage___block_26_v_y;
_q___pip_5160_1_79___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___stage___block_26_v_y : _d___pip_5160_1_79___stage___block_26_v_y;
_q___pip_5160_1_80___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___stage___block_26_v_y : _d___pip_5160_1_80___stage___block_26_v_y;
_q___pip_5160_1_81___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___stage___block_26_v_y : _d___pip_5160_1_81___stage___block_26_v_y;
_q___pip_5160_1_82___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___stage___block_26_v_y : _d___pip_5160_1_82___stage___block_26_v_y;
_q___pip_5160_1_83___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___stage___block_26_v_y : _d___pip_5160_1_83___stage___block_26_v_y;
_q___pip_5160_1_84___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___stage___block_26_v_y : _d___pip_5160_1_84___stage___block_26_v_y;
_q___pip_5160_1_85___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___stage___block_26_v_y : _d___pip_5160_1_85___stage___block_26_v_y;
_q___pip_5160_1_86___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___stage___block_26_v_y : _d___pip_5160_1_86___stage___block_26_v_y;
_q___pip_5160_1_87___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___stage___block_26_v_y : _d___pip_5160_1_87___stage___block_26_v_y;
_q___pip_5160_1_88___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___stage___block_26_v_y : _d___pip_5160_1_88___stage___block_26_v_y;
_q___pip_5160_1_89___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___stage___block_26_v_y : _d___pip_5160_1_89___stage___block_26_v_y;
_q___pip_5160_1_90___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___stage___block_26_v_y : _d___pip_5160_1_90___stage___block_26_v_y;
_q___pip_5160_1_91___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___stage___block_26_v_y : _d___pip_5160_1_91___stage___block_26_v_y;
_q___pip_5160_1_92___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___stage___block_26_v_y : _d___pip_5160_1_92___stage___block_26_v_y;
_q___pip_5160_1_93___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___stage___block_26_v_y : _d___pip_5160_1_93___stage___block_26_v_y;
_q___pip_5160_1_94___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___stage___block_26_v_y : _d___pip_5160_1_94___stage___block_26_v_y;
_q___pip_5160_1_95___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___stage___block_26_v_y : _d___pip_5160_1_95___stage___block_26_v_y;
_q___pip_5160_1_96___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___stage___block_26_v_y : _d___pip_5160_1_96___stage___block_26_v_y;
_q___pip_5160_1_97___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___stage___block_26_v_y : _d___pip_5160_1_97___stage___block_26_v_y;
_q___pip_5160_1_98___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___stage___block_26_v_y : _d___pip_5160_1_98___stage___block_26_v_y;
_q___pip_5160_1_99___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___stage___block_26_v_y : _d___pip_5160_1_99___stage___block_26_v_y;
_q___pip_5160_1_100___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___stage___block_26_v_y : _d___pip_5160_1_100___stage___block_26_v_y;
_q___pip_5160_1_101___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___stage___block_26_v_y : _d___pip_5160_1_101___stage___block_26_v_y;
_q___pip_5160_1_102___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___stage___block_26_v_y : _d___pip_5160_1_102___stage___block_26_v_y;
_q___pip_5160_1_103___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___stage___block_26_v_y : _d___pip_5160_1_103___stage___block_26_v_y;
_q___pip_5160_1_104___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___stage___block_26_v_y : _d___pip_5160_1_104___stage___block_26_v_y;
_q___pip_5160_1_105___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___stage___block_26_v_y : _d___pip_5160_1_105___stage___block_26_v_y;
_q___pip_5160_1_106___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___stage___block_26_v_y : _d___pip_5160_1_106___stage___block_26_v_y;
_q___pip_5160_1_107___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___stage___block_26_v_y : _d___pip_5160_1_107___stage___block_26_v_y;
_q___pip_5160_1_108___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___stage___block_26_v_y : _d___pip_5160_1_108___stage___block_26_v_y;
_q___pip_5160_1_109___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___stage___block_26_v_y : _d___pip_5160_1_109___stage___block_26_v_y;
_q___pip_5160_1_110___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___stage___block_26_v_y : _d___pip_5160_1_110___stage___block_26_v_y;
_q___pip_5160_1_111___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___stage___block_26_v_y : _d___pip_5160_1_111___stage___block_26_v_y;
_q___pip_5160_1_112___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___stage___block_26_v_y : _d___pip_5160_1_112___stage___block_26_v_y;
_q___pip_5160_1_113___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___stage___block_26_v_y : _d___pip_5160_1_113___stage___block_26_v_y;
_q___pip_5160_1_114___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___stage___block_26_v_y : _d___pip_5160_1_114___stage___block_26_v_y;
_q___pip_5160_1_115___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___stage___block_26_v_y : _d___pip_5160_1_115___stage___block_26_v_y;
_q___pip_5160_1_116___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___stage___block_26_v_y : _d___pip_5160_1_116___stage___block_26_v_y;
_q___pip_5160_1_117___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___stage___block_26_v_y : _d___pip_5160_1_117___stage___block_26_v_y;
_q___pip_5160_1_118___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___stage___block_26_v_y : _d___pip_5160_1_118___stage___block_26_v_y;
_q___pip_5160_1_119___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___stage___block_26_v_y : _d___pip_5160_1_119___stage___block_26_v_y;
_q___pip_5160_1_120___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___stage___block_26_v_y : _d___pip_5160_1_120___stage___block_26_v_y;
_q___pip_5160_1_121___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___stage___block_26_v_y : _d___pip_5160_1_121___stage___block_26_v_y;
_q___pip_5160_1_122___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___stage___block_26_v_y : _d___pip_5160_1_122___stage___block_26_v_y;
_q___pip_5160_1_123___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___stage___block_26_v_y : _d___pip_5160_1_123___stage___block_26_v_y;
_q___pip_5160_1_124___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___stage___block_26_v_y : _d___pip_5160_1_124___stage___block_26_v_y;
_q___pip_5160_1_125___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___stage___block_26_v_y : _d___pip_5160_1_125___stage___block_26_v_y;
_q___pip_5160_1_126___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___stage___block_26_v_y : _d___pip_5160_1_126___stage___block_26_v_y;
_q___pip_5160_1_127___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___stage___block_26_v_y : _d___pip_5160_1_127___stage___block_26_v_y;
_q___pip_5160_1_128___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___stage___block_26_v_y : _d___pip_5160_1_128___stage___block_26_v_y;
_q___pip_5160_1_129___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___stage___block_26_v_y : _d___pip_5160_1_129___stage___block_26_v_y;
_q___pip_5160_1_130___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___stage___block_26_v_y : _d___pip_5160_1_130___stage___block_26_v_y;
_q___pip_5160_1_131___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___stage___block_26_v_y : _d___pip_5160_1_131___stage___block_26_v_y;
_q___pip_5160_1_132___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___stage___block_26_v_y : _d___pip_5160_1_132___stage___block_26_v_y;
_q___pip_5160_1_133___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___stage___block_26_v_y : _d___pip_5160_1_133___stage___block_26_v_y;
_q___pip_5160_1_134___stage___block_26_v_y <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___stage___block_26_v_y : _d___pip_5160_1_134___stage___block_26_v_y;
_q___pip_5160_1_4___stage___block_26_v_z <= _d___pip_5160_1_4___stage___block_26_v_z;
_q___pip_5160_1_5___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_26_v_z : _d___pip_5160_1_5___stage___block_26_v_z;
_q___pip_5160_1_6___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_26_v_z : _d___pip_5160_1_6___stage___block_26_v_z;
_q___pip_5160_1_7___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___stage___block_26_v_z : _d___pip_5160_1_7___stage___block_26_v_z;
_q___pip_5160_1_8___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___stage___block_26_v_z : _d___pip_5160_1_8___stage___block_26_v_z;
_q___pip_5160_1_9___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___stage___block_26_v_z : _d___pip_5160_1_9___stage___block_26_v_z;
_q___pip_5160_1_10___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___stage___block_26_v_z : _d___pip_5160_1_10___stage___block_26_v_z;
_q___pip_5160_1_11___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___stage___block_26_v_z : _d___pip_5160_1_11___stage___block_26_v_z;
_q___pip_5160_1_12___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___stage___block_26_v_z : _d___pip_5160_1_12___stage___block_26_v_z;
_q___pip_5160_1_13___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___stage___block_26_v_z : _d___pip_5160_1_13___stage___block_26_v_z;
_q___pip_5160_1_14___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___stage___block_26_v_z : _d___pip_5160_1_14___stage___block_26_v_z;
_q___pip_5160_1_15___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___stage___block_26_v_z : _d___pip_5160_1_15___stage___block_26_v_z;
_q___pip_5160_1_16___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___stage___block_26_v_z : _d___pip_5160_1_16___stage___block_26_v_z;
_q___pip_5160_1_17___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___stage___block_26_v_z : _d___pip_5160_1_17___stage___block_26_v_z;
_q___pip_5160_1_18___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___stage___block_26_v_z : _d___pip_5160_1_18___stage___block_26_v_z;
_q___pip_5160_1_19___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___stage___block_26_v_z : _d___pip_5160_1_19___stage___block_26_v_z;
_q___pip_5160_1_20___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___stage___block_26_v_z : _d___pip_5160_1_20___stage___block_26_v_z;
_q___pip_5160_1_21___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___stage___block_26_v_z : _d___pip_5160_1_21___stage___block_26_v_z;
_q___pip_5160_1_22___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___stage___block_26_v_z : _d___pip_5160_1_22___stage___block_26_v_z;
_q___pip_5160_1_23___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___stage___block_26_v_z : _d___pip_5160_1_23___stage___block_26_v_z;
_q___pip_5160_1_24___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___stage___block_26_v_z : _d___pip_5160_1_24___stage___block_26_v_z;
_q___pip_5160_1_25___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___stage___block_26_v_z : _d___pip_5160_1_25___stage___block_26_v_z;
_q___pip_5160_1_26___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___stage___block_26_v_z : _d___pip_5160_1_26___stage___block_26_v_z;
_q___pip_5160_1_27___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___stage___block_26_v_z : _d___pip_5160_1_27___stage___block_26_v_z;
_q___pip_5160_1_28___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___stage___block_26_v_z : _d___pip_5160_1_28___stage___block_26_v_z;
_q___pip_5160_1_29___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___stage___block_26_v_z : _d___pip_5160_1_29___stage___block_26_v_z;
_q___pip_5160_1_30___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___stage___block_26_v_z : _d___pip_5160_1_30___stage___block_26_v_z;
_q___pip_5160_1_31___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___stage___block_26_v_z : _d___pip_5160_1_31___stage___block_26_v_z;
_q___pip_5160_1_32___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___stage___block_26_v_z : _d___pip_5160_1_32___stage___block_26_v_z;
_q___pip_5160_1_33___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___stage___block_26_v_z : _d___pip_5160_1_33___stage___block_26_v_z;
_q___pip_5160_1_34___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___stage___block_26_v_z : _d___pip_5160_1_34___stage___block_26_v_z;
_q___pip_5160_1_35___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___stage___block_26_v_z : _d___pip_5160_1_35___stage___block_26_v_z;
_q___pip_5160_1_36___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___stage___block_26_v_z : _d___pip_5160_1_36___stage___block_26_v_z;
_q___pip_5160_1_37___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___stage___block_26_v_z : _d___pip_5160_1_37___stage___block_26_v_z;
_q___pip_5160_1_38___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___stage___block_26_v_z : _d___pip_5160_1_38___stage___block_26_v_z;
_q___pip_5160_1_39___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___stage___block_26_v_z : _d___pip_5160_1_39___stage___block_26_v_z;
_q___pip_5160_1_40___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___stage___block_26_v_z : _d___pip_5160_1_40___stage___block_26_v_z;
_q___pip_5160_1_41___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___stage___block_26_v_z : _d___pip_5160_1_41___stage___block_26_v_z;
_q___pip_5160_1_42___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___stage___block_26_v_z : _d___pip_5160_1_42___stage___block_26_v_z;
_q___pip_5160_1_43___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___stage___block_26_v_z : _d___pip_5160_1_43___stage___block_26_v_z;
_q___pip_5160_1_44___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___stage___block_26_v_z : _d___pip_5160_1_44___stage___block_26_v_z;
_q___pip_5160_1_45___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___stage___block_26_v_z : _d___pip_5160_1_45___stage___block_26_v_z;
_q___pip_5160_1_46___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___stage___block_26_v_z : _d___pip_5160_1_46___stage___block_26_v_z;
_q___pip_5160_1_47___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___stage___block_26_v_z : _d___pip_5160_1_47___stage___block_26_v_z;
_q___pip_5160_1_48___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___stage___block_26_v_z : _d___pip_5160_1_48___stage___block_26_v_z;
_q___pip_5160_1_49___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___stage___block_26_v_z : _d___pip_5160_1_49___stage___block_26_v_z;
_q___pip_5160_1_50___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___stage___block_26_v_z : _d___pip_5160_1_50___stage___block_26_v_z;
_q___pip_5160_1_51___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___stage___block_26_v_z : _d___pip_5160_1_51___stage___block_26_v_z;
_q___pip_5160_1_52___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___stage___block_26_v_z : _d___pip_5160_1_52___stage___block_26_v_z;
_q___pip_5160_1_53___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___stage___block_26_v_z : _d___pip_5160_1_53___stage___block_26_v_z;
_q___pip_5160_1_54___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___stage___block_26_v_z : _d___pip_5160_1_54___stage___block_26_v_z;
_q___pip_5160_1_55___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___stage___block_26_v_z : _d___pip_5160_1_55___stage___block_26_v_z;
_q___pip_5160_1_56___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___stage___block_26_v_z : _d___pip_5160_1_56___stage___block_26_v_z;
_q___pip_5160_1_57___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___stage___block_26_v_z : _d___pip_5160_1_57___stage___block_26_v_z;
_q___pip_5160_1_58___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___stage___block_26_v_z : _d___pip_5160_1_58___stage___block_26_v_z;
_q___pip_5160_1_59___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___stage___block_26_v_z : _d___pip_5160_1_59___stage___block_26_v_z;
_q___pip_5160_1_60___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___stage___block_26_v_z : _d___pip_5160_1_60___stage___block_26_v_z;
_q___pip_5160_1_61___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___stage___block_26_v_z : _d___pip_5160_1_61___stage___block_26_v_z;
_q___pip_5160_1_62___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___stage___block_26_v_z : _d___pip_5160_1_62___stage___block_26_v_z;
_q___pip_5160_1_63___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___stage___block_26_v_z : _d___pip_5160_1_63___stage___block_26_v_z;
_q___pip_5160_1_64___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___stage___block_26_v_z : _d___pip_5160_1_64___stage___block_26_v_z;
_q___pip_5160_1_65___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___stage___block_26_v_z : _d___pip_5160_1_65___stage___block_26_v_z;
_q___pip_5160_1_66___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___stage___block_26_v_z : _d___pip_5160_1_66___stage___block_26_v_z;
_q___pip_5160_1_67___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___stage___block_26_v_z : _d___pip_5160_1_67___stage___block_26_v_z;
_q___pip_5160_1_68___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___stage___block_26_v_z : _d___pip_5160_1_68___stage___block_26_v_z;
_q___pip_5160_1_69___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___stage___block_26_v_z : _d___pip_5160_1_69___stage___block_26_v_z;
_q___pip_5160_1_70___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___stage___block_26_v_z : _d___pip_5160_1_70___stage___block_26_v_z;
_q___pip_5160_1_71___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___stage___block_26_v_z : _d___pip_5160_1_71___stage___block_26_v_z;
_q___pip_5160_1_72___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___stage___block_26_v_z : _d___pip_5160_1_72___stage___block_26_v_z;
_q___pip_5160_1_73___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___stage___block_26_v_z : _d___pip_5160_1_73___stage___block_26_v_z;
_q___pip_5160_1_74___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___stage___block_26_v_z : _d___pip_5160_1_74___stage___block_26_v_z;
_q___pip_5160_1_75___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___stage___block_26_v_z : _d___pip_5160_1_75___stage___block_26_v_z;
_q___pip_5160_1_76___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___stage___block_26_v_z : _d___pip_5160_1_76___stage___block_26_v_z;
_q___pip_5160_1_77___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___stage___block_26_v_z : _d___pip_5160_1_77___stage___block_26_v_z;
_q___pip_5160_1_78___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___stage___block_26_v_z : _d___pip_5160_1_78___stage___block_26_v_z;
_q___pip_5160_1_79___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___stage___block_26_v_z : _d___pip_5160_1_79___stage___block_26_v_z;
_q___pip_5160_1_80___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___stage___block_26_v_z : _d___pip_5160_1_80___stage___block_26_v_z;
_q___pip_5160_1_81___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___stage___block_26_v_z : _d___pip_5160_1_81___stage___block_26_v_z;
_q___pip_5160_1_82___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___stage___block_26_v_z : _d___pip_5160_1_82___stage___block_26_v_z;
_q___pip_5160_1_83___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___stage___block_26_v_z : _d___pip_5160_1_83___stage___block_26_v_z;
_q___pip_5160_1_84___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___stage___block_26_v_z : _d___pip_5160_1_84___stage___block_26_v_z;
_q___pip_5160_1_85___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___stage___block_26_v_z : _d___pip_5160_1_85___stage___block_26_v_z;
_q___pip_5160_1_86___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___stage___block_26_v_z : _d___pip_5160_1_86___stage___block_26_v_z;
_q___pip_5160_1_87___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___stage___block_26_v_z : _d___pip_5160_1_87___stage___block_26_v_z;
_q___pip_5160_1_88___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___stage___block_26_v_z : _d___pip_5160_1_88___stage___block_26_v_z;
_q___pip_5160_1_89___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___stage___block_26_v_z : _d___pip_5160_1_89___stage___block_26_v_z;
_q___pip_5160_1_90___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___stage___block_26_v_z : _d___pip_5160_1_90___stage___block_26_v_z;
_q___pip_5160_1_91___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___stage___block_26_v_z : _d___pip_5160_1_91___stage___block_26_v_z;
_q___pip_5160_1_92___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___stage___block_26_v_z : _d___pip_5160_1_92___stage___block_26_v_z;
_q___pip_5160_1_93___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___stage___block_26_v_z : _d___pip_5160_1_93___stage___block_26_v_z;
_q___pip_5160_1_94___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___stage___block_26_v_z : _d___pip_5160_1_94___stage___block_26_v_z;
_q___pip_5160_1_95___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___stage___block_26_v_z : _d___pip_5160_1_95___stage___block_26_v_z;
_q___pip_5160_1_96___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___stage___block_26_v_z : _d___pip_5160_1_96___stage___block_26_v_z;
_q___pip_5160_1_97___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___stage___block_26_v_z : _d___pip_5160_1_97___stage___block_26_v_z;
_q___pip_5160_1_98___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___stage___block_26_v_z : _d___pip_5160_1_98___stage___block_26_v_z;
_q___pip_5160_1_99___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___stage___block_26_v_z : _d___pip_5160_1_99___stage___block_26_v_z;
_q___pip_5160_1_100___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___stage___block_26_v_z : _d___pip_5160_1_100___stage___block_26_v_z;
_q___pip_5160_1_101___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___stage___block_26_v_z : _d___pip_5160_1_101___stage___block_26_v_z;
_q___pip_5160_1_102___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___stage___block_26_v_z : _d___pip_5160_1_102___stage___block_26_v_z;
_q___pip_5160_1_103___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___stage___block_26_v_z : _d___pip_5160_1_103___stage___block_26_v_z;
_q___pip_5160_1_104___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___stage___block_26_v_z : _d___pip_5160_1_104___stage___block_26_v_z;
_q___pip_5160_1_105___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___stage___block_26_v_z : _d___pip_5160_1_105___stage___block_26_v_z;
_q___pip_5160_1_106___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___stage___block_26_v_z : _d___pip_5160_1_106___stage___block_26_v_z;
_q___pip_5160_1_107___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___stage___block_26_v_z : _d___pip_5160_1_107___stage___block_26_v_z;
_q___pip_5160_1_108___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___stage___block_26_v_z : _d___pip_5160_1_108___stage___block_26_v_z;
_q___pip_5160_1_109___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___stage___block_26_v_z : _d___pip_5160_1_109___stage___block_26_v_z;
_q___pip_5160_1_110___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___stage___block_26_v_z : _d___pip_5160_1_110___stage___block_26_v_z;
_q___pip_5160_1_111___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___stage___block_26_v_z : _d___pip_5160_1_111___stage___block_26_v_z;
_q___pip_5160_1_112___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___stage___block_26_v_z : _d___pip_5160_1_112___stage___block_26_v_z;
_q___pip_5160_1_113___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___stage___block_26_v_z : _d___pip_5160_1_113___stage___block_26_v_z;
_q___pip_5160_1_114___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___stage___block_26_v_z : _d___pip_5160_1_114___stage___block_26_v_z;
_q___pip_5160_1_115___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___stage___block_26_v_z : _d___pip_5160_1_115___stage___block_26_v_z;
_q___pip_5160_1_116___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___stage___block_26_v_z : _d___pip_5160_1_116___stage___block_26_v_z;
_q___pip_5160_1_117___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___stage___block_26_v_z : _d___pip_5160_1_117___stage___block_26_v_z;
_q___pip_5160_1_118___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___stage___block_26_v_z : _d___pip_5160_1_118___stage___block_26_v_z;
_q___pip_5160_1_119___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___stage___block_26_v_z : _d___pip_5160_1_119___stage___block_26_v_z;
_q___pip_5160_1_120___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___stage___block_26_v_z : _d___pip_5160_1_120___stage___block_26_v_z;
_q___pip_5160_1_121___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___stage___block_26_v_z : _d___pip_5160_1_121___stage___block_26_v_z;
_q___pip_5160_1_122___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___stage___block_26_v_z : _d___pip_5160_1_122___stage___block_26_v_z;
_q___pip_5160_1_123___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___stage___block_26_v_z : _d___pip_5160_1_123___stage___block_26_v_z;
_q___pip_5160_1_124___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___stage___block_26_v_z : _d___pip_5160_1_124___stage___block_26_v_z;
_q___pip_5160_1_125___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___stage___block_26_v_z : _d___pip_5160_1_125___stage___block_26_v_z;
_q___pip_5160_1_126___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___stage___block_26_v_z : _d___pip_5160_1_126___stage___block_26_v_z;
_q___pip_5160_1_127___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___stage___block_26_v_z : _d___pip_5160_1_127___stage___block_26_v_z;
_q___pip_5160_1_128___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___stage___block_26_v_z : _d___pip_5160_1_128___stage___block_26_v_z;
_q___pip_5160_1_129___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___stage___block_26_v_z : _d___pip_5160_1_129___stage___block_26_v_z;
_q___pip_5160_1_130___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___stage___block_26_v_z : _d___pip_5160_1_130___stage___block_26_v_z;
_q___pip_5160_1_131___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___stage___block_26_v_z : _d___pip_5160_1_131___stage___block_26_v_z;
_q___pip_5160_1_132___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___stage___block_26_v_z : _d___pip_5160_1_132___stage___block_26_v_z;
_q___pip_5160_1_133___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___stage___block_26_v_z : _d___pip_5160_1_133___stage___block_26_v_z;
_q___pip_5160_1_134___stage___block_26_v_z <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___stage___block_26_v_z : _d___pip_5160_1_134___stage___block_26_v_z;
_q___pip_5160_1_0___stage___block_6_clr <= _d___pip_5160_1_0___stage___block_6_clr;
_q___pip_5160_1_1___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_1 == 1 && !_t__stall_fsm___pip_5160_1_1) ? _d___pip_5160_1_0___stage___block_6_clr : _d___pip_5160_1_1___stage___block_6_clr;
_q___pip_5160_1_2___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_2 == 1 && !_t__stall_fsm___pip_5160_1_2) ? _d___pip_5160_1_1___stage___block_6_clr : _d___pip_5160_1_2___stage___block_6_clr;
_q___pip_5160_1_3___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_3 == 1 && !_t__stall_fsm___pip_5160_1_3) ? _d___pip_5160_1_2___stage___block_6_clr : _d___pip_5160_1_3___stage___block_6_clr;
_q___pip_5160_1_4___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_4 == 1 && !_t__stall_fsm___pip_5160_1_4) ? _d___pip_5160_1_3___stage___block_6_clr : _d___pip_5160_1_4___stage___block_6_clr;
_q___pip_5160_1_5___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_6_clr : _d___pip_5160_1_5___stage___block_6_clr;
_q___pip_5160_1_6___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_6_clr : _d___pip_5160_1_6___stage___block_6_clr;
_q___pip_5160_1_7___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___stage___block_6_clr : _d___pip_5160_1_7___stage___block_6_clr;
_q___pip_5160_1_8___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___stage___block_6_clr : _d___pip_5160_1_8___stage___block_6_clr;
_q___pip_5160_1_9___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___stage___block_6_clr : _d___pip_5160_1_9___stage___block_6_clr;
_q___pip_5160_1_10___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___stage___block_6_clr : _d___pip_5160_1_10___stage___block_6_clr;
_q___pip_5160_1_11___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___stage___block_6_clr : _d___pip_5160_1_11___stage___block_6_clr;
_q___pip_5160_1_12___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___stage___block_6_clr : _d___pip_5160_1_12___stage___block_6_clr;
_q___pip_5160_1_13___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___stage___block_6_clr : _d___pip_5160_1_13___stage___block_6_clr;
_q___pip_5160_1_14___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___stage___block_6_clr : _d___pip_5160_1_14___stage___block_6_clr;
_q___pip_5160_1_15___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___stage___block_6_clr : _d___pip_5160_1_15___stage___block_6_clr;
_q___pip_5160_1_16___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___stage___block_6_clr : _d___pip_5160_1_16___stage___block_6_clr;
_q___pip_5160_1_17___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___stage___block_6_clr : _d___pip_5160_1_17___stage___block_6_clr;
_q___pip_5160_1_18___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___stage___block_6_clr : _d___pip_5160_1_18___stage___block_6_clr;
_q___pip_5160_1_19___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___stage___block_6_clr : _d___pip_5160_1_19___stage___block_6_clr;
_q___pip_5160_1_20___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___stage___block_6_clr : _d___pip_5160_1_20___stage___block_6_clr;
_q___pip_5160_1_21___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___stage___block_6_clr : _d___pip_5160_1_21___stage___block_6_clr;
_q___pip_5160_1_22___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___stage___block_6_clr : _d___pip_5160_1_22___stage___block_6_clr;
_q___pip_5160_1_23___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___stage___block_6_clr : _d___pip_5160_1_23___stage___block_6_clr;
_q___pip_5160_1_24___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___stage___block_6_clr : _d___pip_5160_1_24___stage___block_6_clr;
_q___pip_5160_1_25___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___stage___block_6_clr : _d___pip_5160_1_25___stage___block_6_clr;
_q___pip_5160_1_26___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___stage___block_6_clr : _d___pip_5160_1_26___stage___block_6_clr;
_q___pip_5160_1_27___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___stage___block_6_clr : _d___pip_5160_1_27___stage___block_6_clr;
_q___pip_5160_1_28___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___stage___block_6_clr : _d___pip_5160_1_28___stage___block_6_clr;
_q___pip_5160_1_29___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___stage___block_6_clr : _d___pip_5160_1_29___stage___block_6_clr;
_q___pip_5160_1_30___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___stage___block_6_clr : _d___pip_5160_1_30___stage___block_6_clr;
_q___pip_5160_1_31___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___stage___block_6_clr : _d___pip_5160_1_31___stage___block_6_clr;
_q___pip_5160_1_32___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___stage___block_6_clr : _d___pip_5160_1_32___stage___block_6_clr;
_q___pip_5160_1_33___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___stage___block_6_clr : _d___pip_5160_1_33___stage___block_6_clr;
_q___pip_5160_1_34___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___stage___block_6_clr : _d___pip_5160_1_34___stage___block_6_clr;
_q___pip_5160_1_35___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___stage___block_6_clr : _d___pip_5160_1_35___stage___block_6_clr;
_q___pip_5160_1_36___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___stage___block_6_clr : _d___pip_5160_1_36___stage___block_6_clr;
_q___pip_5160_1_37___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___stage___block_6_clr : _d___pip_5160_1_37___stage___block_6_clr;
_q___pip_5160_1_38___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___stage___block_6_clr : _d___pip_5160_1_38___stage___block_6_clr;
_q___pip_5160_1_39___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___stage___block_6_clr : _d___pip_5160_1_39___stage___block_6_clr;
_q___pip_5160_1_40___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___stage___block_6_clr : _d___pip_5160_1_40___stage___block_6_clr;
_q___pip_5160_1_41___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___stage___block_6_clr : _d___pip_5160_1_41___stage___block_6_clr;
_q___pip_5160_1_42___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___stage___block_6_clr : _d___pip_5160_1_42___stage___block_6_clr;
_q___pip_5160_1_43___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___stage___block_6_clr : _d___pip_5160_1_43___stage___block_6_clr;
_q___pip_5160_1_44___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___stage___block_6_clr : _d___pip_5160_1_44___stage___block_6_clr;
_q___pip_5160_1_45___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___stage___block_6_clr : _d___pip_5160_1_45___stage___block_6_clr;
_q___pip_5160_1_46___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___stage___block_6_clr : _d___pip_5160_1_46___stage___block_6_clr;
_q___pip_5160_1_47___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___stage___block_6_clr : _d___pip_5160_1_47___stage___block_6_clr;
_q___pip_5160_1_48___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___stage___block_6_clr : _d___pip_5160_1_48___stage___block_6_clr;
_q___pip_5160_1_49___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___stage___block_6_clr : _d___pip_5160_1_49___stage___block_6_clr;
_q___pip_5160_1_50___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___stage___block_6_clr : _d___pip_5160_1_50___stage___block_6_clr;
_q___pip_5160_1_51___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___stage___block_6_clr : _d___pip_5160_1_51___stage___block_6_clr;
_q___pip_5160_1_52___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___stage___block_6_clr : _d___pip_5160_1_52___stage___block_6_clr;
_q___pip_5160_1_53___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___stage___block_6_clr : _d___pip_5160_1_53___stage___block_6_clr;
_q___pip_5160_1_54___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___stage___block_6_clr : _d___pip_5160_1_54___stage___block_6_clr;
_q___pip_5160_1_55___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___stage___block_6_clr : _d___pip_5160_1_55___stage___block_6_clr;
_q___pip_5160_1_56___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___stage___block_6_clr : _d___pip_5160_1_56___stage___block_6_clr;
_q___pip_5160_1_57___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___stage___block_6_clr : _d___pip_5160_1_57___stage___block_6_clr;
_q___pip_5160_1_58___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___stage___block_6_clr : _d___pip_5160_1_58___stage___block_6_clr;
_q___pip_5160_1_59___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___stage___block_6_clr : _d___pip_5160_1_59___stage___block_6_clr;
_q___pip_5160_1_60___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___stage___block_6_clr : _d___pip_5160_1_60___stage___block_6_clr;
_q___pip_5160_1_61___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___stage___block_6_clr : _d___pip_5160_1_61___stage___block_6_clr;
_q___pip_5160_1_62___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___stage___block_6_clr : _d___pip_5160_1_62___stage___block_6_clr;
_q___pip_5160_1_63___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___stage___block_6_clr : _d___pip_5160_1_63___stage___block_6_clr;
_q___pip_5160_1_64___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___stage___block_6_clr : _d___pip_5160_1_64___stage___block_6_clr;
_q___pip_5160_1_65___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___stage___block_6_clr : _d___pip_5160_1_65___stage___block_6_clr;
_q___pip_5160_1_66___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___stage___block_6_clr : _d___pip_5160_1_66___stage___block_6_clr;
_q___pip_5160_1_67___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___stage___block_6_clr : _d___pip_5160_1_67___stage___block_6_clr;
_q___pip_5160_1_68___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___stage___block_6_clr : _d___pip_5160_1_68___stage___block_6_clr;
_q___pip_5160_1_69___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___stage___block_6_clr : _d___pip_5160_1_69___stage___block_6_clr;
_q___pip_5160_1_70___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___stage___block_6_clr : _d___pip_5160_1_70___stage___block_6_clr;
_q___pip_5160_1_71___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___stage___block_6_clr : _d___pip_5160_1_71___stage___block_6_clr;
_q___pip_5160_1_72___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___stage___block_6_clr : _d___pip_5160_1_72___stage___block_6_clr;
_q___pip_5160_1_73___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___stage___block_6_clr : _d___pip_5160_1_73___stage___block_6_clr;
_q___pip_5160_1_74___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___stage___block_6_clr : _d___pip_5160_1_74___stage___block_6_clr;
_q___pip_5160_1_75___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___stage___block_6_clr : _d___pip_5160_1_75___stage___block_6_clr;
_q___pip_5160_1_76___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___stage___block_6_clr : _d___pip_5160_1_76___stage___block_6_clr;
_q___pip_5160_1_77___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___stage___block_6_clr : _d___pip_5160_1_77___stage___block_6_clr;
_q___pip_5160_1_78___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___stage___block_6_clr : _d___pip_5160_1_78___stage___block_6_clr;
_q___pip_5160_1_79___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___stage___block_6_clr : _d___pip_5160_1_79___stage___block_6_clr;
_q___pip_5160_1_80___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___stage___block_6_clr : _d___pip_5160_1_80___stage___block_6_clr;
_q___pip_5160_1_81___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___stage___block_6_clr : _d___pip_5160_1_81___stage___block_6_clr;
_q___pip_5160_1_82___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___stage___block_6_clr : _d___pip_5160_1_82___stage___block_6_clr;
_q___pip_5160_1_83___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___stage___block_6_clr : _d___pip_5160_1_83___stage___block_6_clr;
_q___pip_5160_1_84___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___stage___block_6_clr : _d___pip_5160_1_84___stage___block_6_clr;
_q___pip_5160_1_85___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___stage___block_6_clr : _d___pip_5160_1_85___stage___block_6_clr;
_q___pip_5160_1_86___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___stage___block_6_clr : _d___pip_5160_1_86___stage___block_6_clr;
_q___pip_5160_1_87___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___stage___block_6_clr : _d___pip_5160_1_87___stage___block_6_clr;
_q___pip_5160_1_88___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___stage___block_6_clr : _d___pip_5160_1_88___stage___block_6_clr;
_q___pip_5160_1_89___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___stage___block_6_clr : _d___pip_5160_1_89___stage___block_6_clr;
_q___pip_5160_1_90___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___stage___block_6_clr : _d___pip_5160_1_90___stage___block_6_clr;
_q___pip_5160_1_91___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___stage___block_6_clr : _d___pip_5160_1_91___stage___block_6_clr;
_q___pip_5160_1_92___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___stage___block_6_clr : _d___pip_5160_1_92___stage___block_6_clr;
_q___pip_5160_1_93___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___stage___block_6_clr : _d___pip_5160_1_93___stage___block_6_clr;
_q___pip_5160_1_94___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___stage___block_6_clr : _d___pip_5160_1_94___stage___block_6_clr;
_q___pip_5160_1_95___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___stage___block_6_clr : _d___pip_5160_1_95___stage___block_6_clr;
_q___pip_5160_1_96___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___stage___block_6_clr : _d___pip_5160_1_96___stage___block_6_clr;
_q___pip_5160_1_97___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___stage___block_6_clr : _d___pip_5160_1_97___stage___block_6_clr;
_q___pip_5160_1_98___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___stage___block_6_clr : _d___pip_5160_1_98___stage___block_6_clr;
_q___pip_5160_1_99___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___stage___block_6_clr : _d___pip_5160_1_99___stage___block_6_clr;
_q___pip_5160_1_100___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___stage___block_6_clr : _d___pip_5160_1_100___stage___block_6_clr;
_q___pip_5160_1_101___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___stage___block_6_clr : _d___pip_5160_1_101___stage___block_6_clr;
_q___pip_5160_1_102___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___stage___block_6_clr : _d___pip_5160_1_102___stage___block_6_clr;
_q___pip_5160_1_103___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___stage___block_6_clr : _d___pip_5160_1_103___stage___block_6_clr;
_q___pip_5160_1_104___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___stage___block_6_clr : _d___pip_5160_1_104___stage___block_6_clr;
_q___pip_5160_1_105___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___stage___block_6_clr : _d___pip_5160_1_105___stage___block_6_clr;
_q___pip_5160_1_106___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___stage___block_6_clr : _d___pip_5160_1_106___stage___block_6_clr;
_q___pip_5160_1_107___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___stage___block_6_clr : _d___pip_5160_1_107___stage___block_6_clr;
_q___pip_5160_1_108___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___stage___block_6_clr : _d___pip_5160_1_108___stage___block_6_clr;
_q___pip_5160_1_109___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___stage___block_6_clr : _d___pip_5160_1_109___stage___block_6_clr;
_q___pip_5160_1_110___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___stage___block_6_clr : _d___pip_5160_1_110___stage___block_6_clr;
_q___pip_5160_1_111___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___stage___block_6_clr : _d___pip_5160_1_111___stage___block_6_clr;
_q___pip_5160_1_112___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___stage___block_6_clr : _d___pip_5160_1_112___stage___block_6_clr;
_q___pip_5160_1_113___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___stage___block_6_clr : _d___pip_5160_1_113___stage___block_6_clr;
_q___pip_5160_1_114___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___stage___block_6_clr : _d___pip_5160_1_114___stage___block_6_clr;
_q___pip_5160_1_115___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___stage___block_6_clr : _d___pip_5160_1_115___stage___block_6_clr;
_q___pip_5160_1_116___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___stage___block_6_clr : _d___pip_5160_1_116___stage___block_6_clr;
_q___pip_5160_1_117___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___stage___block_6_clr : _d___pip_5160_1_117___stage___block_6_clr;
_q___pip_5160_1_118___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___stage___block_6_clr : _d___pip_5160_1_118___stage___block_6_clr;
_q___pip_5160_1_119___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___stage___block_6_clr : _d___pip_5160_1_119___stage___block_6_clr;
_q___pip_5160_1_120___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___stage___block_6_clr : _d___pip_5160_1_120___stage___block_6_clr;
_q___pip_5160_1_121___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___stage___block_6_clr : _d___pip_5160_1_121___stage___block_6_clr;
_q___pip_5160_1_122___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___stage___block_6_clr : _d___pip_5160_1_122___stage___block_6_clr;
_q___pip_5160_1_123___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___stage___block_6_clr : _d___pip_5160_1_123___stage___block_6_clr;
_q___pip_5160_1_124___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___stage___block_6_clr : _d___pip_5160_1_124___stage___block_6_clr;
_q___pip_5160_1_125___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___stage___block_6_clr : _d___pip_5160_1_125___stage___block_6_clr;
_q___pip_5160_1_126___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___stage___block_6_clr : _d___pip_5160_1_126___stage___block_6_clr;
_q___pip_5160_1_127___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___stage___block_6_clr : _d___pip_5160_1_127___stage___block_6_clr;
_q___pip_5160_1_128___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___stage___block_6_clr : _d___pip_5160_1_128___stage___block_6_clr;
_q___pip_5160_1_129___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___stage___block_6_clr : _d___pip_5160_1_129___stage___block_6_clr;
_q___pip_5160_1_130___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___stage___block_6_clr : _d___pip_5160_1_130___stage___block_6_clr;
_q___pip_5160_1_131___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___stage___block_6_clr : _d___pip_5160_1_131___stage___block_6_clr;
_q___pip_5160_1_132___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___stage___block_6_clr : _d___pip_5160_1_132___stage___block_6_clr;
_q___pip_5160_1_133___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___stage___block_6_clr : _d___pip_5160_1_133___stage___block_6_clr;
_q___pip_5160_1_134___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___stage___block_6_clr : _d___pip_5160_1_134___stage___block_6_clr;
_q___pip_5160_1_135___stage___block_6_clr <= (_d__idx_fsm___pip_5160_1_135 == 1 && !_t__stall_fsm___pip_5160_1_135) ? _d___pip_5160_1_134___stage___block_6_clr : _d___pip_5160_1_135___stage___block_6_clr;
_q___pip_5160_1_0___stage___block_6_dist <= _d___pip_5160_1_0___stage___block_6_dist;
_q___pip_5160_1_1___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_1 == 1 && !_t__stall_fsm___pip_5160_1_1) ? _d___pip_5160_1_0___stage___block_6_dist : _d___pip_5160_1_1___stage___block_6_dist;
_q___pip_5160_1_2___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_2 == 1 && !_t__stall_fsm___pip_5160_1_2) ? _d___pip_5160_1_1___stage___block_6_dist : _d___pip_5160_1_2___stage___block_6_dist;
_q___pip_5160_1_3___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_3 == 1 && !_t__stall_fsm___pip_5160_1_3) ? _d___pip_5160_1_2___stage___block_6_dist : _d___pip_5160_1_3___stage___block_6_dist;
_q___pip_5160_1_4___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_4 == 1 && !_t__stall_fsm___pip_5160_1_4) ? _d___pip_5160_1_3___stage___block_6_dist : _d___pip_5160_1_4___stage___block_6_dist;
_q___pip_5160_1_5___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_6_dist : _d___pip_5160_1_5___stage___block_6_dist;
_q___pip_5160_1_6___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_6_dist : _d___pip_5160_1_6___stage___block_6_dist;
_q___pip_5160_1_7___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___stage___block_6_dist : _d___pip_5160_1_7___stage___block_6_dist;
_q___pip_5160_1_8___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___stage___block_6_dist : _d___pip_5160_1_8___stage___block_6_dist;
_q___pip_5160_1_9___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___stage___block_6_dist : _d___pip_5160_1_9___stage___block_6_dist;
_q___pip_5160_1_10___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___stage___block_6_dist : _d___pip_5160_1_10___stage___block_6_dist;
_q___pip_5160_1_11___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___stage___block_6_dist : _d___pip_5160_1_11___stage___block_6_dist;
_q___pip_5160_1_12___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___stage___block_6_dist : _d___pip_5160_1_12___stage___block_6_dist;
_q___pip_5160_1_13___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___stage___block_6_dist : _d___pip_5160_1_13___stage___block_6_dist;
_q___pip_5160_1_14___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___stage___block_6_dist : _d___pip_5160_1_14___stage___block_6_dist;
_q___pip_5160_1_15___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___stage___block_6_dist : _d___pip_5160_1_15___stage___block_6_dist;
_q___pip_5160_1_16___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___stage___block_6_dist : _d___pip_5160_1_16___stage___block_6_dist;
_q___pip_5160_1_17___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___stage___block_6_dist : _d___pip_5160_1_17___stage___block_6_dist;
_q___pip_5160_1_18___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___stage___block_6_dist : _d___pip_5160_1_18___stage___block_6_dist;
_q___pip_5160_1_19___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___stage___block_6_dist : _d___pip_5160_1_19___stage___block_6_dist;
_q___pip_5160_1_20___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___stage___block_6_dist : _d___pip_5160_1_20___stage___block_6_dist;
_q___pip_5160_1_21___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___stage___block_6_dist : _d___pip_5160_1_21___stage___block_6_dist;
_q___pip_5160_1_22___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___stage___block_6_dist : _d___pip_5160_1_22___stage___block_6_dist;
_q___pip_5160_1_23___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___stage___block_6_dist : _d___pip_5160_1_23___stage___block_6_dist;
_q___pip_5160_1_24___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___stage___block_6_dist : _d___pip_5160_1_24___stage___block_6_dist;
_q___pip_5160_1_25___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___stage___block_6_dist : _d___pip_5160_1_25___stage___block_6_dist;
_q___pip_5160_1_26___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___stage___block_6_dist : _d___pip_5160_1_26___stage___block_6_dist;
_q___pip_5160_1_27___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___stage___block_6_dist : _d___pip_5160_1_27___stage___block_6_dist;
_q___pip_5160_1_28___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___stage___block_6_dist : _d___pip_5160_1_28___stage___block_6_dist;
_q___pip_5160_1_29___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___stage___block_6_dist : _d___pip_5160_1_29___stage___block_6_dist;
_q___pip_5160_1_30___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___stage___block_6_dist : _d___pip_5160_1_30___stage___block_6_dist;
_q___pip_5160_1_31___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___stage___block_6_dist : _d___pip_5160_1_31___stage___block_6_dist;
_q___pip_5160_1_32___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___stage___block_6_dist : _d___pip_5160_1_32___stage___block_6_dist;
_q___pip_5160_1_33___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___stage___block_6_dist : _d___pip_5160_1_33___stage___block_6_dist;
_q___pip_5160_1_34___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___stage___block_6_dist : _d___pip_5160_1_34___stage___block_6_dist;
_q___pip_5160_1_35___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___stage___block_6_dist : _d___pip_5160_1_35___stage___block_6_dist;
_q___pip_5160_1_36___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___stage___block_6_dist : _d___pip_5160_1_36___stage___block_6_dist;
_q___pip_5160_1_37___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___stage___block_6_dist : _d___pip_5160_1_37___stage___block_6_dist;
_q___pip_5160_1_38___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___stage___block_6_dist : _d___pip_5160_1_38___stage___block_6_dist;
_q___pip_5160_1_39___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___stage___block_6_dist : _d___pip_5160_1_39___stage___block_6_dist;
_q___pip_5160_1_40___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___stage___block_6_dist : _d___pip_5160_1_40___stage___block_6_dist;
_q___pip_5160_1_41___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___stage___block_6_dist : _d___pip_5160_1_41___stage___block_6_dist;
_q___pip_5160_1_42___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___stage___block_6_dist : _d___pip_5160_1_42___stage___block_6_dist;
_q___pip_5160_1_43___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___stage___block_6_dist : _d___pip_5160_1_43___stage___block_6_dist;
_q___pip_5160_1_44___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___stage___block_6_dist : _d___pip_5160_1_44___stage___block_6_dist;
_q___pip_5160_1_45___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___stage___block_6_dist : _d___pip_5160_1_45___stage___block_6_dist;
_q___pip_5160_1_46___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___stage___block_6_dist : _d___pip_5160_1_46___stage___block_6_dist;
_q___pip_5160_1_47___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___stage___block_6_dist : _d___pip_5160_1_47___stage___block_6_dist;
_q___pip_5160_1_48___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___stage___block_6_dist : _d___pip_5160_1_48___stage___block_6_dist;
_q___pip_5160_1_49___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___stage___block_6_dist : _d___pip_5160_1_49___stage___block_6_dist;
_q___pip_5160_1_50___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___stage___block_6_dist : _d___pip_5160_1_50___stage___block_6_dist;
_q___pip_5160_1_51___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___stage___block_6_dist : _d___pip_5160_1_51___stage___block_6_dist;
_q___pip_5160_1_52___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___stage___block_6_dist : _d___pip_5160_1_52___stage___block_6_dist;
_q___pip_5160_1_53___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___stage___block_6_dist : _d___pip_5160_1_53___stage___block_6_dist;
_q___pip_5160_1_54___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___stage___block_6_dist : _d___pip_5160_1_54___stage___block_6_dist;
_q___pip_5160_1_55___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___stage___block_6_dist : _d___pip_5160_1_55___stage___block_6_dist;
_q___pip_5160_1_56___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___stage___block_6_dist : _d___pip_5160_1_56___stage___block_6_dist;
_q___pip_5160_1_57___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___stage___block_6_dist : _d___pip_5160_1_57___stage___block_6_dist;
_q___pip_5160_1_58___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___stage___block_6_dist : _d___pip_5160_1_58___stage___block_6_dist;
_q___pip_5160_1_59___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___stage___block_6_dist : _d___pip_5160_1_59___stage___block_6_dist;
_q___pip_5160_1_60___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___stage___block_6_dist : _d___pip_5160_1_60___stage___block_6_dist;
_q___pip_5160_1_61___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___stage___block_6_dist : _d___pip_5160_1_61___stage___block_6_dist;
_q___pip_5160_1_62___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___stage___block_6_dist : _d___pip_5160_1_62___stage___block_6_dist;
_q___pip_5160_1_63___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___stage___block_6_dist : _d___pip_5160_1_63___stage___block_6_dist;
_q___pip_5160_1_64___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___stage___block_6_dist : _d___pip_5160_1_64___stage___block_6_dist;
_q___pip_5160_1_65___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___stage___block_6_dist : _d___pip_5160_1_65___stage___block_6_dist;
_q___pip_5160_1_66___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___stage___block_6_dist : _d___pip_5160_1_66___stage___block_6_dist;
_q___pip_5160_1_67___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___stage___block_6_dist : _d___pip_5160_1_67___stage___block_6_dist;
_q___pip_5160_1_68___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___stage___block_6_dist : _d___pip_5160_1_68___stage___block_6_dist;
_q___pip_5160_1_69___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___stage___block_6_dist : _d___pip_5160_1_69___stage___block_6_dist;
_q___pip_5160_1_70___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___stage___block_6_dist : _d___pip_5160_1_70___stage___block_6_dist;
_q___pip_5160_1_71___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___stage___block_6_dist : _d___pip_5160_1_71___stage___block_6_dist;
_q___pip_5160_1_72___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___stage___block_6_dist : _d___pip_5160_1_72___stage___block_6_dist;
_q___pip_5160_1_73___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___stage___block_6_dist : _d___pip_5160_1_73___stage___block_6_dist;
_q___pip_5160_1_74___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___stage___block_6_dist : _d___pip_5160_1_74___stage___block_6_dist;
_q___pip_5160_1_75___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___stage___block_6_dist : _d___pip_5160_1_75___stage___block_6_dist;
_q___pip_5160_1_76___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___stage___block_6_dist : _d___pip_5160_1_76___stage___block_6_dist;
_q___pip_5160_1_77___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___stage___block_6_dist : _d___pip_5160_1_77___stage___block_6_dist;
_q___pip_5160_1_78___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___stage___block_6_dist : _d___pip_5160_1_78___stage___block_6_dist;
_q___pip_5160_1_79___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___stage___block_6_dist : _d___pip_5160_1_79___stage___block_6_dist;
_q___pip_5160_1_80___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___stage___block_6_dist : _d___pip_5160_1_80___stage___block_6_dist;
_q___pip_5160_1_81___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___stage___block_6_dist : _d___pip_5160_1_81___stage___block_6_dist;
_q___pip_5160_1_82___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___stage___block_6_dist : _d___pip_5160_1_82___stage___block_6_dist;
_q___pip_5160_1_83___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___stage___block_6_dist : _d___pip_5160_1_83___stage___block_6_dist;
_q___pip_5160_1_84___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___stage___block_6_dist : _d___pip_5160_1_84___stage___block_6_dist;
_q___pip_5160_1_85___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___stage___block_6_dist : _d___pip_5160_1_85___stage___block_6_dist;
_q___pip_5160_1_86___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___stage___block_6_dist : _d___pip_5160_1_86___stage___block_6_dist;
_q___pip_5160_1_87___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___stage___block_6_dist : _d___pip_5160_1_87___stage___block_6_dist;
_q___pip_5160_1_88___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___stage___block_6_dist : _d___pip_5160_1_88___stage___block_6_dist;
_q___pip_5160_1_89___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___stage___block_6_dist : _d___pip_5160_1_89___stage___block_6_dist;
_q___pip_5160_1_90___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___stage___block_6_dist : _d___pip_5160_1_90___stage___block_6_dist;
_q___pip_5160_1_91___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___stage___block_6_dist : _d___pip_5160_1_91___stage___block_6_dist;
_q___pip_5160_1_92___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___stage___block_6_dist : _d___pip_5160_1_92___stage___block_6_dist;
_q___pip_5160_1_93___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___stage___block_6_dist : _d___pip_5160_1_93___stage___block_6_dist;
_q___pip_5160_1_94___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___stage___block_6_dist : _d___pip_5160_1_94___stage___block_6_dist;
_q___pip_5160_1_95___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___stage___block_6_dist : _d___pip_5160_1_95___stage___block_6_dist;
_q___pip_5160_1_96___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___stage___block_6_dist : _d___pip_5160_1_96___stage___block_6_dist;
_q___pip_5160_1_97___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___stage___block_6_dist : _d___pip_5160_1_97___stage___block_6_dist;
_q___pip_5160_1_98___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___stage___block_6_dist : _d___pip_5160_1_98___stage___block_6_dist;
_q___pip_5160_1_99___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___stage___block_6_dist : _d___pip_5160_1_99___stage___block_6_dist;
_q___pip_5160_1_100___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___stage___block_6_dist : _d___pip_5160_1_100___stage___block_6_dist;
_q___pip_5160_1_101___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___stage___block_6_dist : _d___pip_5160_1_101___stage___block_6_dist;
_q___pip_5160_1_102___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___stage___block_6_dist : _d___pip_5160_1_102___stage___block_6_dist;
_q___pip_5160_1_103___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___stage___block_6_dist : _d___pip_5160_1_103___stage___block_6_dist;
_q___pip_5160_1_104___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___stage___block_6_dist : _d___pip_5160_1_104___stage___block_6_dist;
_q___pip_5160_1_105___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___stage___block_6_dist : _d___pip_5160_1_105___stage___block_6_dist;
_q___pip_5160_1_106___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___stage___block_6_dist : _d___pip_5160_1_106___stage___block_6_dist;
_q___pip_5160_1_107___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___stage___block_6_dist : _d___pip_5160_1_107___stage___block_6_dist;
_q___pip_5160_1_108___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___stage___block_6_dist : _d___pip_5160_1_108___stage___block_6_dist;
_q___pip_5160_1_109___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___stage___block_6_dist : _d___pip_5160_1_109___stage___block_6_dist;
_q___pip_5160_1_110___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___stage___block_6_dist : _d___pip_5160_1_110___stage___block_6_dist;
_q___pip_5160_1_111___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___stage___block_6_dist : _d___pip_5160_1_111___stage___block_6_dist;
_q___pip_5160_1_112___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___stage___block_6_dist : _d___pip_5160_1_112___stage___block_6_dist;
_q___pip_5160_1_113___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___stage___block_6_dist : _d___pip_5160_1_113___stage___block_6_dist;
_q___pip_5160_1_114___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___stage___block_6_dist : _d___pip_5160_1_114___stage___block_6_dist;
_q___pip_5160_1_115___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___stage___block_6_dist : _d___pip_5160_1_115___stage___block_6_dist;
_q___pip_5160_1_116___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___stage___block_6_dist : _d___pip_5160_1_116___stage___block_6_dist;
_q___pip_5160_1_117___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___stage___block_6_dist : _d___pip_5160_1_117___stage___block_6_dist;
_q___pip_5160_1_118___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___stage___block_6_dist : _d___pip_5160_1_118___stage___block_6_dist;
_q___pip_5160_1_119___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___stage___block_6_dist : _d___pip_5160_1_119___stage___block_6_dist;
_q___pip_5160_1_120___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___stage___block_6_dist : _d___pip_5160_1_120___stage___block_6_dist;
_q___pip_5160_1_121___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___stage___block_6_dist : _d___pip_5160_1_121___stage___block_6_dist;
_q___pip_5160_1_122___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___stage___block_6_dist : _d___pip_5160_1_122___stage___block_6_dist;
_q___pip_5160_1_123___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___stage___block_6_dist : _d___pip_5160_1_123___stage___block_6_dist;
_q___pip_5160_1_124___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___stage___block_6_dist : _d___pip_5160_1_124___stage___block_6_dist;
_q___pip_5160_1_125___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___stage___block_6_dist : _d___pip_5160_1_125___stage___block_6_dist;
_q___pip_5160_1_126___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___stage___block_6_dist : _d___pip_5160_1_126___stage___block_6_dist;
_q___pip_5160_1_127___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___stage___block_6_dist : _d___pip_5160_1_127___stage___block_6_dist;
_q___pip_5160_1_128___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___stage___block_6_dist : _d___pip_5160_1_128___stage___block_6_dist;
_q___pip_5160_1_129___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___stage___block_6_dist : _d___pip_5160_1_129___stage___block_6_dist;
_q___pip_5160_1_130___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___stage___block_6_dist : _d___pip_5160_1_130___stage___block_6_dist;
_q___pip_5160_1_131___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___stage___block_6_dist : _d___pip_5160_1_131___stage___block_6_dist;
_q___pip_5160_1_132___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___stage___block_6_dist : _d___pip_5160_1_132___stage___block_6_dist;
_q___pip_5160_1_133___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___stage___block_6_dist : _d___pip_5160_1_133___stage___block_6_dist;
_q___pip_5160_1_134___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___stage___block_6_dist : _d___pip_5160_1_134___stage___block_6_dist;
_q___pip_5160_1_135___stage___block_6_dist <= (_d__idx_fsm___pip_5160_1_135 == 1 && !_t__stall_fsm___pip_5160_1_135) ? _d___pip_5160_1_134___stage___block_6_dist : _d___pip_5160_1_135___stage___block_6_dist;
_q___pip_5160_1_0___stage___block_6_inside <= _d___pip_5160_1_0___stage___block_6_inside;
_q___pip_5160_1_1___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_1 == 1 && !_t__stall_fsm___pip_5160_1_1) ? _d___pip_5160_1_0___stage___block_6_inside : _d___pip_5160_1_1___stage___block_6_inside;
_q___pip_5160_1_2___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_2 == 1 && !_t__stall_fsm___pip_5160_1_2) ? _d___pip_5160_1_1___stage___block_6_inside : _d___pip_5160_1_2___stage___block_6_inside;
_q___pip_5160_1_3___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_3 == 1 && !_t__stall_fsm___pip_5160_1_3) ? _d___pip_5160_1_2___stage___block_6_inside : _d___pip_5160_1_3___stage___block_6_inside;
_q___pip_5160_1_4___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_4 == 1 && !_t__stall_fsm___pip_5160_1_4) ? _d___pip_5160_1_3___stage___block_6_inside : _d___pip_5160_1_4___stage___block_6_inside;
_q___pip_5160_1_5___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_6_inside : _d___pip_5160_1_5___stage___block_6_inside;
_q___pip_5160_1_6___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_6_inside : _d___pip_5160_1_6___stage___block_6_inside;
_q___pip_5160_1_7___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_7 == 1 && !_t__stall_fsm___pip_5160_1_7) ? _d___pip_5160_1_6___stage___block_6_inside : _d___pip_5160_1_7___stage___block_6_inside;
_q___pip_5160_1_8___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_8 == 1 && !_t__stall_fsm___pip_5160_1_8) ? _d___pip_5160_1_7___stage___block_6_inside : _d___pip_5160_1_8___stage___block_6_inside;
_q___pip_5160_1_9___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_9 == 1 && !_t__stall_fsm___pip_5160_1_9) ? _d___pip_5160_1_8___stage___block_6_inside : _d___pip_5160_1_9___stage___block_6_inside;
_q___pip_5160_1_10___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_10 == 1 && !_t__stall_fsm___pip_5160_1_10) ? _d___pip_5160_1_9___stage___block_6_inside : _d___pip_5160_1_10___stage___block_6_inside;
_q___pip_5160_1_11___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_11 == 1 && !_t__stall_fsm___pip_5160_1_11) ? _d___pip_5160_1_10___stage___block_6_inside : _d___pip_5160_1_11___stage___block_6_inside;
_q___pip_5160_1_12___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_12 == 1 && !_t__stall_fsm___pip_5160_1_12) ? _d___pip_5160_1_11___stage___block_6_inside : _d___pip_5160_1_12___stage___block_6_inside;
_q___pip_5160_1_13___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_13 == 1 && !_t__stall_fsm___pip_5160_1_13) ? _d___pip_5160_1_12___stage___block_6_inside : _d___pip_5160_1_13___stage___block_6_inside;
_q___pip_5160_1_14___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_14 == 1 && !_t__stall_fsm___pip_5160_1_14) ? _d___pip_5160_1_13___stage___block_6_inside : _d___pip_5160_1_14___stage___block_6_inside;
_q___pip_5160_1_15___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_15 == 1 && !_t__stall_fsm___pip_5160_1_15) ? _d___pip_5160_1_14___stage___block_6_inside : _d___pip_5160_1_15___stage___block_6_inside;
_q___pip_5160_1_16___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_16 == 1 && !_t__stall_fsm___pip_5160_1_16) ? _d___pip_5160_1_15___stage___block_6_inside : _d___pip_5160_1_16___stage___block_6_inside;
_q___pip_5160_1_17___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_17 == 1 && !_t__stall_fsm___pip_5160_1_17) ? _d___pip_5160_1_16___stage___block_6_inside : _d___pip_5160_1_17___stage___block_6_inside;
_q___pip_5160_1_18___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_18 == 1 && !_t__stall_fsm___pip_5160_1_18) ? _d___pip_5160_1_17___stage___block_6_inside : _d___pip_5160_1_18___stage___block_6_inside;
_q___pip_5160_1_19___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_19 == 1 && !_t__stall_fsm___pip_5160_1_19) ? _d___pip_5160_1_18___stage___block_6_inside : _d___pip_5160_1_19___stage___block_6_inside;
_q___pip_5160_1_20___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_20 == 1 && !_t__stall_fsm___pip_5160_1_20) ? _d___pip_5160_1_19___stage___block_6_inside : _d___pip_5160_1_20___stage___block_6_inside;
_q___pip_5160_1_21___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_21 == 1 && !_t__stall_fsm___pip_5160_1_21) ? _d___pip_5160_1_20___stage___block_6_inside : _d___pip_5160_1_21___stage___block_6_inside;
_q___pip_5160_1_22___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_22 == 1 && !_t__stall_fsm___pip_5160_1_22) ? _d___pip_5160_1_21___stage___block_6_inside : _d___pip_5160_1_22___stage___block_6_inside;
_q___pip_5160_1_23___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_23 == 1 && !_t__stall_fsm___pip_5160_1_23) ? _d___pip_5160_1_22___stage___block_6_inside : _d___pip_5160_1_23___stage___block_6_inside;
_q___pip_5160_1_24___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_24 == 1 && !_t__stall_fsm___pip_5160_1_24) ? _d___pip_5160_1_23___stage___block_6_inside : _d___pip_5160_1_24___stage___block_6_inside;
_q___pip_5160_1_25___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_25 == 1 && !_t__stall_fsm___pip_5160_1_25) ? _d___pip_5160_1_24___stage___block_6_inside : _d___pip_5160_1_25___stage___block_6_inside;
_q___pip_5160_1_26___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_26 == 1 && !_t__stall_fsm___pip_5160_1_26) ? _d___pip_5160_1_25___stage___block_6_inside : _d___pip_5160_1_26___stage___block_6_inside;
_q___pip_5160_1_27___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_27 == 1 && !_t__stall_fsm___pip_5160_1_27) ? _d___pip_5160_1_26___stage___block_6_inside : _d___pip_5160_1_27___stage___block_6_inside;
_q___pip_5160_1_28___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_28 == 1 && !_t__stall_fsm___pip_5160_1_28) ? _d___pip_5160_1_27___stage___block_6_inside : _d___pip_5160_1_28___stage___block_6_inside;
_q___pip_5160_1_29___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_29 == 1 && !_t__stall_fsm___pip_5160_1_29) ? _d___pip_5160_1_28___stage___block_6_inside : _d___pip_5160_1_29___stage___block_6_inside;
_q___pip_5160_1_30___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_30 == 1 && !_t__stall_fsm___pip_5160_1_30) ? _d___pip_5160_1_29___stage___block_6_inside : _d___pip_5160_1_30___stage___block_6_inside;
_q___pip_5160_1_31___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_31 == 1 && !_t__stall_fsm___pip_5160_1_31) ? _d___pip_5160_1_30___stage___block_6_inside : _d___pip_5160_1_31___stage___block_6_inside;
_q___pip_5160_1_32___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_32 == 1 && !_t__stall_fsm___pip_5160_1_32) ? _d___pip_5160_1_31___stage___block_6_inside : _d___pip_5160_1_32___stage___block_6_inside;
_q___pip_5160_1_33___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_33 == 1 && !_t__stall_fsm___pip_5160_1_33) ? _d___pip_5160_1_32___stage___block_6_inside : _d___pip_5160_1_33___stage___block_6_inside;
_q___pip_5160_1_34___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_34 == 1 && !_t__stall_fsm___pip_5160_1_34) ? _d___pip_5160_1_33___stage___block_6_inside : _d___pip_5160_1_34___stage___block_6_inside;
_q___pip_5160_1_35___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_35 == 1 && !_t__stall_fsm___pip_5160_1_35) ? _d___pip_5160_1_34___stage___block_6_inside : _d___pip_5160_1_35___stage___block_6_inside;
_q___pip_5160_1_36___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_36 == 1 && !_t__stall_fsm___pip_5160_1_36) ? _d___pip_5160_1_35___stage___block_6_inside : _d___pip_5160_1_36___stage___block_6_inside;
_q___pip_5160_1_37___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_37 == 1 && !_t__stall_fsm___pip_5160_1_37) ? _d___pip_5160_1_36___stage___block_6_inside : _d___pip_5160_1_37___stage___block_6_inside;
_q___pip_5160_1_38___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_38 == 1 && !_t__stall_fsm___pip_5160_1_38) ? _d___pip_5160_1_37___stage___block_6_inside : _d___pip_5160_1_38___stage___block_6_inside;
_q___pip_5160_1_39___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_39 == 1 && !_t__stall_fsm___pip_5160_1_39) ? _d___pip_5160_1_38___stage___block_6_inside : _d___pip_5160_1_39___stage___block_6_inside;
_q___pip_5160_1_40___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_40 == 1 && !_t__stall_fsm___pip_5160_1_40) ? _d___pip_5160_1_39___stage___block_6_inside : _d___pip_5160_1_40___stage___block_6_inside;
_q___pip_5160_1_41___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_41 == 1 && !_t__stall_fsm___pip_5160_1_41) ? _d___pip_5160_1_40___stage___block_6_inside : _d___pip_5160_1_41___stage___block_6_inside;
_q___pip_5160_1_42___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_42 == 1 && !_t__stall_fsm___pip_5160_1_42) ? _d___pip_5160_1_41___stage___block_6_inside : _d___pip_5160_1_42___stage___block_6_inside;
_q___pip_5160_1_43___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_43 == 1 && !_t__stall_fsm___pip_5160_1_43) ? _d___pip_5160_1_42___stage___block_6_inside : _d___pip_5160_1_43___stage___block_6_inside;
_q___pip_5160_1_44___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_44 == 1 && !_t__stall_fsm___pip_5160_1_44) ? _d___pip_5160_1_43___stage___block_6_inside : _d___pip_5160_1_44___stage___block_6_inside;
_q___pip_5160_1_45___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_45 == 1 && !_t__stall_fsm___pip_5160_1_45) ? _d___pip_5160_1_44___stage___block_6_inside : _d___pip_5160_1_45___stage___block_6_inside;
_q___pip_5160_1_46___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_46 == 1 && !_t__stall_fsm___pip_5160_1_46) ? _d___pip_5160_1_45___stage___block_6_inside : _d___pip_5160_1_46___stage___block_6_inside;
_q___pip_5160_1_47___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_47 == 1 && !_t__stall_fsm___pip_5160_1_47) ? _d___pip_5160_1_46___stage___block_6_inside : _d___pip_5160_1_47___stage___block_6_inside;
_q___pip_5160_1_48___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_48 == 1 && !_t__stall_fsm___pip_5160_1_48) ? _d___pip_5160_1_47___stage___block_6_inside : _d___pip_5160_1_48___stage___block_6_inside;
_q___pip_5160_1_49___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_49 == 1 && !_t__stall_fsm___pip_5160_1_49) ? _d___pip_5160_1_48___stage___block_6_inside : _d___pip_5160_1_49___stage___block_6_inside;
_q___pip_5160_1_50___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_50 == 1 && !_t__stall_fsm___pip_5160_1_50) ? _d___pip_5160_1_49___stage___block_6_inside : _d___pip_5160_1_50___stage___block_6_inside;
_q___pip_5160_1_51___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_51 == 1 && !_t__stall_fsm___pip_5160_1_51) ? _d___pip_5160_1_50___stage___block_6_inside : _d___pip_5160_1_51___stage___block_6_inside;
_q___pip_5160_1_52___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_52 == 1 && !_t__stall_fsm___pip_5160_1_52) ? _d___pip_5160_1_51___stage___block_6_inside : _d___pip_5160_1_52___stage___block_6_inside;
_q___pip_5160_1_53___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_53 == 1 && !_t__stall_fsm___pip_5160_1_53) ? _d___pip_5160_1_52___stage___block_6_inside : _d___pip_5160_1_53___stage___block_6_inside;
_q___pip_5160_1_54___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_54 == 1 && !_t__stall_fsm___pip_5160_1_54) ? _d___pip_5160_1_53___stage___block_6_inside : _d___pip_5160_1_54___stage___block_6_inside;
_q___pip_5160_1_55___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_55 == 1 && !_t__stall_fsm___pip_5160_1_55) ? _d___pip_5160_1_54___stage___block_6_inside : _d___pip_5160_1_55___stage___block_6_inside;
_q___pip_5160_1_56___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_56 == 1 && !_t__stall_fsm___pip_5160_1_56) ? _d___pip_5160_1_55___stage___block_6_inside : _d___pip_5160_1_56___stage___block_6_inside;
_q___pip_5160_1_57___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_57 == 1 && !_t__stall_fsm___pip_5160_1_57) ? _d___pip_5160_1_56___stage___block_6_inside : _d___pip_5160_1_57___stage___block_6_inside;
_q___pip_5160_1_58___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_58 == 1 && !_t__stall_fsm___pip_5160_1_58) ? _d___pip_5160_1_57___stage___block_6_inside : _d___pip_5160_1_58___stage___block_6_inside;
_q___pip_5160_1_59___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_59 == 1 && !_t__stall_fsm___pip_5160_1_59) ? _d___pip_5160_1_58___stage___block_6_inside : _d___pip_5160_1_59___stage___block_6_inside;
_q___pip_5160_1_60___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_60 == 1 && !_t__stall_fsm___pip_5160_1_60) ? _d___pip_5160_1_59___stage___block_6_inside : _d___pip_5160_1_60___stage___block_6_inside;
_q___pip_5160_1_61___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_61 == 1 && !_t__stall_fsm___pip_5160_1_61) ? _d___pip_5160_1_60___stage___block_6_inside : _d___pip_5160_1_61___stage___block_6_inside;
_q___pip_5160_1_62___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_62 == 1 && !_t__stall_fsm___pip_5160_1_62) ? _d___pip_5160_1_61___stage___block_6_inside : _d___pip_5160_1_62___stage___block_6_inside;
_q___pip_5160_1_63___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_63 == 1 && !_t__stall_fsm___pip_5160_1_63) ? _d___pip_5160_1_62___stage___block_6_inside : _d___pip_5160_1_63___stage___block_6_inside;
_q___pip_5160_1_64___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_64 == 1 && !_t__stall_fsm___pip_5160_1_64) ? _d___pip_5160_1_63___stage___block_6_inside : _d___pip_5160_1_64___stage___block_6_inside;
_q___pip_5160_1_65___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_65 == 1 && !_t__stall_fsm___pip_5160_1_65) ? _d___pip_5160_1_64___stage___block_6_inside : _d___pip_5160_1_65___stage___block_6_inside;
_q___pip_5160_1_66___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_66 == 1 && !_t__stall_fsm___pip_5160_1_66) ? _d___pip_5160_1_65___stage___block_6_inside : _d___pip_5160_1_66___stage___block_6_inside;
_q___pip_5160_1_67___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_67 == 1 && !_t__stall_fsm___pip_5160_1_67) ? _d___pip_5160_1_66___stage___block_6_inside : _d___pip_5160_1_67___stage___block_6_inside;
_q___pip_5160_1_68___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_68 == 1 && !_t__stall_fsm___pip_5160_1_68) ? _d___pip_5160_1_67___stage___block_6_inside : _d___pip_5160_1_68___stage___block_6_inside;
_q___pip_5160_1_69___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_69 == 1 && !_t__stall_fsm___pip_5160_1_69) ? _d___pip_5160_1_68___stage___block_6_inside : _d___pip_5160_1_69___stage___block_6_inside;
_q___pip_5160_1_70___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_70 == 1 && !_t__stall_fsm___pip_5160_1_70) ? _d___pip_5160_1_69___stage___block_6_inside : _d___pip_5160_1_70___stage___block_6_inside;
_q___pip_5160_1_71___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_71 == 1 && !_t__stall_fsm___pip_5160_1_71) ? _d___pip_5160_1_70___stage___block_6_inside : _d___pip_5160_1_71___stage___block_6_inside;
_q___pip_5160_1_72___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_72 == 1 && !_t__stall_fsm___pip_5160_1_72) ? _d___pip_5160_1_71___stage___block_6_inside : _d___pip_5160_1_72___stage___block_6_inside;
_q___pip_5160_1_73___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_73 == 1 && !_t__stall_fsm___pip_5160_1_73) ? _d___pip_5160_1_72___stage___block_6_inside : _d___pip_5160_1_73___stage___block_6_inside;
_q___pip_5160_1_74___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_74 == 1 && !_t__stall_fsm___pip_5160_1_74) ? _d___pip_5160_1_73___stage___block_6_inside : _d___pip_5160_1_74___stage___block_6_inside;
_q___pip_5160_1_75___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_75 == 1 && !_t__stall_fsm___pip_5160_1_75) ? _d___pip_5160_1_74___stage___block_6_inside : _d___pip_5160_1_75___stage___block_6_inside;
_q___pip_5160_1_76___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_76 == 1 && !_t__stall_fsm___pip_5160_1_76) ? _d___pip_5160_1_75___stage___block_6_inside : _d___pip_5160_1_76___stage___block_6_inside;
_q___pip_5160_1_77___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_77 == 1 && !_t__stall_fsm___pip_5160_1_77) ? _d___pip_5160_1_76___stage___block_6_inside : _d___pip_5160_1_77___stage___block_6_inside;
_q___pip_5160_1_78___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_78 == 1 && !_t__stall_fsm___pip_5160_1_78) ? _d___pip_5160_1_77___stage___block_6_inside : _d___pip_5160_1_78___stage___block_6_inside;
_q___pip_5160_1_79___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_79 == 1 && !_t__stall_fsm___pip_5160_1_79) ? _d___pip_5160_1_78___stage___block_6_inside : _d___pip_5160_1_79___stage___block_6_inside;
_q___pip_5160_1_80___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_80 == 1 && !_t__stall_fsm___pip_5160_1_80) ? _d___pip_5160_1_79___stage___block_6_inside : _d___pip_5160_1_80___stage___block_6_inside;
_q___pip_5160_1_81___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_81 == 1 && !_t__stall_fsm___pip_5160_1_81) ? _d___pip_5160_1_80___stage___block_6_inside : _d___pip_5160_1_81___stage___block_6_inside;
_q___pip_5160_1_82___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_82 == 1 && !_t__stall_fsm___pip_5160_1_82) ? _d___pip_5160_1_81___stage___block_6_inside : _d___pip_5160_1_82___stage___block_6_inside;
_q___pip_5160_1_83___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_83 == 1 && !_t__stall_fsm___pip_5160_1_83) ? _d___pip_5160_1_82___stage___block_6_inside : _d___pip_5160_1_83___stage___block_6_inside;
_q___pip_5160_1_84___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_84 == 1 && !_t__stall_fsm___pip_5160_1_84) ? _d___pip_5160_1_83___stage___block_6_inside : _d___pip_5160_1_84___stage___block_6_inside;
_q___pip_5160_1_85___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_85 == 1 && !_t__stall_fsm___pip_5160_1_85) ? _d___pip_5160_1_84___stage___block_6_inside : _d___pip_5160_1_85___stage___block_6_inside;
_q___pip_5160_1_86___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_86 == 1 && !_t__stall_fsm___pip_5160_1_86) ? _d___pip_5160_1_85___stage___block_6_inside : _d___pip_5160_1_86___stage___block_6_inside;
_q___pip_5160_1_87___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_87 == 1 && !_t__stall_fsm___pip_5160_1_87) ? _d___pip_5160_1_86___stage___block_6_inside : _d___pip_5160_1_87___stage___block_6_inside;
_q___pip_5160_1_88___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_88 == 1 && !_t__stall_fsm___pip_5160_1_88) ? _d___pip_5160_1_87___stage___block_6_inside : _d___pip_5160_1_88___stage___block_6_inside;
_q___pip_5160_1_89___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_89 == 1 && !_t__stall_fsm___pip_5160_1_89) ? _d___pip_5160_1_88___stage___block_6_inside : _d___pip_5160_1_89___stage___block_6_inside;
_q___pip_5160_1_90___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_90 == 1 && !_t__stall_fsm___pip_5160_1_90) ? _d___pip_5160_1_89___stage___block_6_inside : _d___pip_5160_1_90___stage___block_6_inside;
_q___pip_5160_1_91___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_91 == 1 && !_t__stall_fsm___pip_5160_1_91) ? _d___pip_5160_1_90___stage___block_6_inside : _d___pip_5160_1_91___stage___block_6_inside;
_q___pip_5160_1_92___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_92 == 1 && !_t__stall_fsm___pip_5160_1_92) ? _d___pip_5160_1_91___stage___block_6_inside : _d___pip_5160_1_92___stage___block_6_inside;
_q___pip_5160_1_93___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_93 == 1 && !_t__stall_fsm___pip_5160_1_93) ? _d___pip_5160_1_92___stage___block_6_inside : _d___pip_5160_1_93___stage___block_6_inside;
_q___pip_5160_1_94___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_94 == 1 && !_t__stall_fsm___pip_5160_1_94) ? _d___pip_5160_1_93___stage___block_6_inside : _d___pip_5160_1_94___stage___block_6_inside;
_q___pip_5160_1_95___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_95 == 1 && !_t__stall_fsm___pip_5160_1_95) ? _d___pip_5160_1_94___stage___block_6_inside : _d___pip_5160_1_95___stage___block_6_inside;
_q___pip_5160_1_96___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_96 == 1 && !_t__stall_fsm___pip_5160_1_96) ? _d___pip_5160_1_95___stage___block_6_inside : _d___pip_5160_1_96___stage___block_6_inside;
_q___pip_5160_1_97___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_97 == 1 && !_t__stall_fsm___pip_5160_1_97) ? _d___pip_5160_1_96___stage___block_6_inside : _d___pip_5160_1_97___stage___block_6_inside;
_q___pip_5160_1_98___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_98 == 1 && !_t__stall_fsm___pip_5160_1_98) ? _d___pip_5160_1_97___stage___block_6_inside : _d___pip_5160_1_98___stage___block_6_inside;
_q___pip_5160_1_99___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_99 == 1 && !_t__stall_fsm___pip_5160_1_99) ? _d___pip_5160_1_98___stage___block_6_inside : _d___pip_5160_1_99___stage___block_6_inside;
_q___pip_5160_1_100___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_100 == 1 && !_t__stall_fsm___pip_5160_1_100) ? _d___pip_5160_1_99___stage___block_6_inside : _d___pip_5160_1_100___stage___block_6_inside;
_q___pip_5160_1_101___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_101 == 1 && !_t__stall_fsm___pip_5160_1_101) ? _d___pip_5160_1_100___stage___block_6_inside : _d___pip_5160_1_101___stage___block_6_inside;
_q___pip_5160_1_102___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_102 == 1 && !_t__stall_fsm___pip_5160_1_102) ? _d___pip_5160_1_101___stage___block_6_inside : _d___pip_5160_1_102___stage___block_6_inside;
_q___pip_5160_1_103___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_103 == 1 && !_t__stall_fsm___pip_5160_1_103) ? _d___pip_5160_1_102___stage___block_6_inside : _d___pip_5160_1_103___stage___block_6_inside;
_q___pip_5160_1_104___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_104 == 1 && !_t__stall_fsm___pip_5160_1_104) ? _d___pip_5160_1_103___stage___block_6_inside : _d___pip_5160_1_104___stage___block_6_inside;
_q___pip_5160_1_105___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_105 == 1 && !_t__stall_fsm___pip_5160_1_105) ? _d___pip_5160_1_104___stage___block_6_inside : _d___pip_5160_1_105___stage___block_6_inside;
_q___pip_5160_1_106___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_106 == 1 && !_t__stall_fsm___pip_5160_1_106) ? _d___pip_5160_1_105___stage___block_6_inside : _d___pip_5160_1_106___stage___block_6_inside;
_q___pip_5160_1_107___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_107 == 1 && !_t__stall_fsm___pip_5160_1_107) ? _d___pip_5160_1_106___stage___block_6_inside : _d___pip_5160_1_107___stage___block_6_inside;
_q___pip_5160_1_108___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_108 == 1 && !_t__stall_fsm___pip_5160_1_108) ? _d___pip_5160_1_107___stage___block_6_inside : _d___pip_5160_1_108___stage___block_6_inside;
_q___pip_5160_1_109___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_109 == 1 && !_t__stall_fsm___pip_5160_1_109) ? _d___pip_5160_1_108___stage___block_6_inside : _d___pip_5160_1_109___stage___block_6_inside;
_q___pip_5160_1_110___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_110 == 1 && !_t__stall_fsm___pip_5160_1_110) ? _d___pip_5160_1_109___stage___block_6_inside : _d___pip_5160_1_110___stage___block_6_inside;
_q___pip_5160_1_111___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_111 == 1 && !_t__stall_fsm___pip_5160_1_111) ? _d___pip_5160_1_110___stage___block_6_inside : _d___pip_5160_1_111___stage___block_6_inside;
_q___pip_5160_1_112___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_112 == 1 && !_t__stall_fsm___pip_5160_1_112) ? _d___pip_5160_1_111___stage___block_6_inside : _d___pip_5160_1_112___stage___block_6_inside;
_q___pip_5160_1_113___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_113 == 1 && !_t__stall_fsm___pip_5160_1_113) ? _d___pip_5160_1_112___stage___block_6_inside : _d___pip_5160_1_113___stage___block_6_inside;
_q___pip_5160_1_114___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_114 == 1 && !_t__stall_fsm___pip_5160_1_114) ? _d___pip_5160_1_113___stage___block_6_inside : _d___pip_5160_1_114___stage___block_6_inside;
_q___pip_5160_1_115___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_115 == 1 && !_t__stall_fsm___pip_5160_1_115) ? _d___pip_5160_1_114___stage___block_6_inside : _d___pip_5160_1_115___stage___block_6_inside;
_q___pip_5160_1_116___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_116 == 1 && !_t__stall_fsm___pip_5160_1_116) ? _d___pip_5160_1_115___stage___block_6_inside : _d___pip_5160_1_116___stage___block_6_inside;
_q___pip_5160_1_117___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_117 == 1 && !_t__stall_fsm___pip_5160_1_117) ? _d___pip_5160_1_116___stage___block_6_inside : _d___pip_5160_1_117___stage___block_6_inside;
_q___pip_5160_1_118___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_118 == 1 && !_t__stall_fsm___pip_5160_1_118) ? _d___pip_5160_1_117___stage___block_6_inside : _d___pip_5160_1_118___stage___block_6_inside;
_q___pip_5160_1_119___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_119 == 1 && !_t__stall_fsm___pip_5160_1_119) ? _d___pip_5160_1_118___stage___block_6_inside : _d___pip_5160_1_119___stage___block_6_inside;
_q___pip_5160_1_120___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_120 == 1 && !_t__stall_fsm___pip_5160_1_120) ? _d___pip_5160_1_119___stage___block_6_inside : _d___pip_5160_1_120___stage___block_6_inside;
_q___pip_5160_1_121___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_121 == 1 && !_t__stall_fsm___pip_5160_1_121) ? _d___pip_5160_1_120___stage___block_6_inside : _d___pip_5160_1_121___stage___block_6_inside;
_q___pip_5160_1_122___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_122 == 1 && !_t__stall_fsm___pip_5160_1_122) ? _d___pip_5160_1_121___stage___block_6_inside : _d___pip_5160_1_122___stage___block_6_inside;
_q___pip_5160_1_123___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_123 == 1 && !_t__stall_fsm___pip_5160_1_123) ? _d___pip_5160_1_122___stage___block_6_inside : _d___pip_5160_1_123___stage___block_6_inside;
_q___pip_5160_1_124___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_124 == 1 && !_t__stall_fsm___pip_5160_1_124) ? _d___pip_5160_1_123___stage___block_6_inside : _d___pip_5160_1_124___stage___block_6_inside;
_q___pip_5160_1_125___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_125 == 1 && !_t__stall_fsm___pip_5160_1_125) ? _d___pip_5160_1_124___stage___block_6_inside : _d___pip_5160_1_125___stage___block_6_inside;
_q___pip_5160_1_126___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_126 == 1 && !_t__stall_fsm___pip_5160_1_126) ? _d___pip_5160_1_125___stage___block_6_inside : _d___pip_5160_1_126___stage___block_6_inside;
_q___pip_5160_1_127___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_127 == 1 && !_t__stall_fsm___pip_5160_1_127) ? _d___pip_5160_1_126___stage___block_6_inside : _d___pip_5160_1_127___stage___block_6_inside;
_q___pip_5160_1_128___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_128 == 1 && !_t__stall_fsm___pip_5160_1_128) ? _d___pip_5160_1_127___stage___block_6_inside : _d___pip_5160_1_128___stage___block_6_inside;
_q___pip_5160_1_129___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_129 == 1 && !_t__stall_fsm___pip_5160_1_129) ? _d___pip_5160_1_128___stage___block_6_inside : _d___pip_5160_1_129___stage___block_6_inside;
_q___pip_5160_1_130___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_130 == 1 && !_t__stall_fsm___pip_5160_1_130) ? _d___pip_5160_1_129___stage___block_6_inside : _d___pip_5160_1_130___stage___block_6_inside;
_q___pip_5160_1_131___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_131 == 1 && !_t__stall_fsm___pip_5160_1_131) ? _d___pip_5160_1_130___stage___block_6_inside : _d___pip_5160_1_131___stage___block_6_inside;
_q___pip_5160_1_132___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_132 == 1 && !_t__stall_fsm___pip_5160_1_132) ? _d___pip_5160_1_131___stage___block_6_inside : _d___pip_5160_1_132___stage___block_6_inside;
_q___pip_5160_1_133___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_133 == 1 && !_t__stall_fsm___pip_5160_1_133) ? _d___pip_5160_1_132___stage___block_6_inside : _d___pip_5160_1_133___stage___block_6_inside;
_q___pip_5160_1_134___stage___block_6_inside <= (_d__idx_fsm___pip_5160_1_134 == 1 && !_t__stall_fsm___pip_5160_1_134) ? _d___pip_5160_1_133___stage___block_6_inside : _d___pip_5160_1_134___stage___block_6_inside;
_q___pip_5160_1_0___stage___block_6_view_x <= _d___pip_5160_1_0___stage___block_6_view_x;
_q___pip_5160_1_1___stage___block_6_view_x <= (_d__idx_fsm___pip_5160_1_1 == 1 && !_t__stall_fsm___pip_5160_1_1) ? _d___pip_5160_1_0___stage___block_6_view_x : _d___pip_5160_1_1___stage___block_6_view_x;
_q___pip_5160_1_2___stage___block_6_view_x <= (_d__idx_fsm___pip_5160_1_2 == 1 && !_t__stall_fsm___pip_5160_1_2) ? _d___pip_5160_1_1___stage___block_6_view_x : _d___pip_5160_1_2___stage___block_6_view_x;
_q___pip_5160_1_3___stage___block_6_view_x <= (_d__idx_fsm___pip_5160_1_3 == 1 && !_t__stall_fsm___pip_5160_1_3) ? _d___pip_5160_1_2___stage___block_6_view_x : _d___pip_5160_1_3___stage___block_6_view_x;
_q___pip_5160_1_0___stage___block_6_view_y <= _d___pip_5160_1_0___stage___block_6_view_y;
_q___pip_5160_1_1___stage___block_6_view_y <= (_d__idx_fsm___pip_5160_1_1 == 1 && !_t__stall_fsm___pip_5160_1_1) ? _d___pip_5160_1_0___stage___block_6_view_y : _d___pip_5160_1_1___stage___block_6_view_y;
_q___pip_5160_1_2___stage___block_6_view_y <= (_d__idx_fsm___pip_5160_1_2 == 1 && !_t__stall_fsm___pip_5160_1_2) ? _d___pip_5160_1_1___stage___block_6_view_y : _d___pip_5160_1_2___stage___block_6_view_y;
_q___pip_5160_1_3___stage___block_6_view_y <= (_d__idx_fsm___pip_5160_1_3 == 1 && !_t__stall_fsm___pip_5160_1_3) ? _d___pip_5160_1_2___stage___block_6_view_y : _d___pip_5160_1_3___stage___block_6_view_y;
_q___pip_5160_1_4___stage___block_6_view_y <= (_d__idx_fsm___pip_5160_1_4 == 1 && !_t__stall_fsm___pip_5160_1_4) ? _d___pip_5160_1_3___stage___block_6_view_y : _d___pip_5160_1_4___stage___block_6_view_y;
_q___pip_5160_1_0___stage___block_6_view_z <= _d___pip_5160_1_0___stage___block_6_view_z;
_q___pip_5160_1_1___stage___block_6_view_z <= (_d__idx_fsm___pip_5160_1_1 == 1 && !_t__stall_fsm___pip_5160_1_1) ? _d___pip_5160_1_0___stage___block_6_view_z : _d___pip_5160_1_1___stage___block_6_view_z;
_q___pip_5160_1_2___stage___block_6_view_z <= (_d__idx_fsm___pip_5160_1_2 == 1 && !_t__stall_fsm___pip_5160_1_2) ? _d___pip_5160_1_1___stage___block_6_view_z : _d___pip_5160_1_2___stage___block_6_view_z;
_q___pip_5160_1_3___stage___block_6_view_z <= (_d__idx_fsm___pip_5160_1_3 == 1 && !_t__stall_fsm___pip_5160_1_3) ? _d___pip_5160_1_2___stage___block_6_view_z : _d___pip_5160_1_3___stage___block_6_view_z;
_q___pip_5160_1_0___stage___block_6_vxsz <= _d___pip_5160_1_0___stage___block_6_vxsz;
_q___pip_5160_1_1___stage___block_6_vxsz <= (_d__idx_fsm___pip_5160_1_1 == 1 && !_t__stall_fsm___pip_5160_1_1) ? _d___pip_5160_1_0___stage___block_6_vxsz : _d___pip_5160_1_1___stage___block_6_vxsz;
_q___pip_5160_1_2___stage___block_6_vxsz <= (_d__idx_fsm___pip_5160_1_2 == 1 && !_t__stall_fsm___pip_5160_1_2) ? _d___pip_5160_1_1___stage___block_6_vxsz : _d___pip_5160_1_2___stage___block_6_vxsz;
_q___pip_5160_1_3___stage___block_6_vxsz <= (_d__idx_fsm___pip_5160_1_3 == 1 && !_t__stall_fsm___pip_5160_1_3) ? _d___pip_5160_1_2___stage___block_6_vxsz : _d___pip_5160_1_3___stage___block_6_vxsz;
_q___pip_5160_1_4___stage___block_6_vxsz <= (_d__idx_fsm___pip_5160_1_4 == 1 && !_t__stall_fsm___pip_5160_1_4) ? _d___pip_5160_1_3___stage___block_6_vxsz : _d___pip_5160_1_4___stage___block_6_vxsz;
_q___pip_5160_1_5___stage___block_6_vxsz <= (_d__idx_fsm___pip_5160_1_5 == 1 && !_t__stall_fsm___pip_5160_1_5) ? _d___pip_5160_1_4___stage___block_6_vxsz : _d___pip_5160_1_5___stage___block_6_vxsz;
_q___pip_5160_1_6___stage___block_6_vxsz <= (_d__idx_fsm___pip_5160_1_6 == 1 && !_t__stall_fsm___pip_5160_1_6) ? _d___pip_5160_1_5___stage___block_6_vxsz : _d___pip_5160_1_6___stage___block_6_vxsz;
_q___pip_5160_1_1___stage___block_7_cs0 <= _d___pip_5160_1_1___stage___block_7_cs0;
_q___pip_5160_1_2___stage___block_7_cs0 <= (_d__idx_fsm___pip_5160_1_2 == 1 && !_t__stall_fsm___pip_5160_1_2) ? _d___pip_5160_1_1___stage___block_7_cs0 : _d___pip_5160_1_2___stage___block_7_cs0;
_q___pip_5160_1_3___stage___block_7_cs0 <= (_d__idx_fsm___pip_5160_1_3 == 1 && !_t__stall_fsm___pip_5160_1_3) ? _d___pip_5160_1_2___stage___block_7_cs0 : _d___pip_5160_1_3___stage___block_7_cs0;
_q___pip_5160_1_1___stage___block_7_ss0 <= _d___pip_5160_1_1___stage___block_7_ss0;
_q___pip_5160_1_2___stage___block_7_ss0 <= (_d__idx_fsm___pip_5160_1_2 == 1 && !_t__stall_fsm___pip_5160_1_2) ? _d___pip_5160_1_1___stage___block_7_ss0 : _d___pip_5160_1_2___stage___block_7_ss0;
_q___pip_5160_1_3___stage___block_7_ss0 <= (_d__idx_fsm___pip_5160_1_3 == 1 && !_t__stall_fsm___pip_5160_1_3) ? _d___pip_5160_1_2___stage___block_7_ss0 : _d___pip_5160_1_3___stage___block_7_ss0;
_q_pix_r <= _d_pix_r;
_q_pix_g <= _d_pix_g;
_q_pix_b <= _d_pix_b;
_q__idx_fsm0 <= reset ? 0 : ( ~_autorun ? 1 : _d__idx_fsm0);
_autorun <= reset ? 0 : 1;
_q__idx_fsm___pip_5160_1_0 <= reset ? 0 : _d__idx_fsm___pip_5160_1_0;
_q__full_fsm___pip_5160_1_0 <= reset ? 0 : _d__full_fsm___pip_5160_1_0;
_q__idx_fsm___pip_5160_1_1 <= reset ? 0 : _d__idx_fsm___pip_5160_1_1;
_q__full_fsm___pip_5160_1_1 <= reset ? 0 : _d__full_fsm___pip_5160_1_1;
_q__idx_fsm___pip_5160_1_2 <= reset ? 0 : _d__idx_fsm___pip_5160_1_2;
_q__full_fsm___pip_5160_1_2 <= reset ? 0 : _d__full_fsm___pip_5160_1_2;
_q__idx_fsm___pip_5160_1_3 <= reset ? 0 : _d__idx_fsm___pip_5160_1_3;
_q__full_fsm___pip_5160_1_3 <= reset ? 0 : _d__full_fsm___pip_5160_1_3;
_q__idx_fsm___pip_5160_1_4 <= reset ? 0 : _d__idx_fsm___pip_5160_1_4;
_q__full_fsm___pip_5160_1_4 <= reset ? 0 : _d__full_fsm___pip_5160_1_4;
_q__idx_fsm___pip_5160_1_5 <= reset ? 0 : _d__idx_fsm___pip_5160_1_5;
_q__full_fsm___pip_5160_1_5 <= reset ? 0 : _d__full_fsm___pip_5160_1_5;
_q__idx_fsm___pip_5160_1_6 <= reset ? 0 : _d__idx_fsm___pip_5160_1_6;
_q__full_fsm___pip_5160_1_6 <= reset ? 0 : _d__full_fsm___pip_5160_1_6;
_q__idx_fsm___pip_5160_1_7 <= reset ? 0 : _d__idx_fsm___pip_5160_1_7;
_q__full_fsm___pip_5160_1_7 <= reset ? 0 : _d__full_fsm___pip_5160_1_7;
_q__idx_fsm___pip_5160_1_8 <= reset ? 0 : _d__idx_fsm___pip_5160_1_8;
_q__full_fsm___pip_5160_1_8 <= reset ? 0 : _d__full_fsm___pip_5160_1_8;
_q__idx_fsm___pip_5160_1_9 <= reset ? 0 : _d__idx_fsm___pip_5160_1_9;
_q__full_fsm___pip_5160_1_9 <= reset ? 0 : _d__full_fsm___pip_5160_1_9;
_q__idx_fsm___pip_5160_1_10 <= reset ? 0 : _d__idx_fsm___pip_5160_1_10;
_q__full_fsm___pip_5160_1_10 <= reset ? 0 : _d__full_fsm___pip_5160_1_10;
_q__idx_fsm___pip_5160_1_11 <= reset ? 0 : _d__idx_fsm___pip_5160_1_11;
_q__full_fsm___pip_5160_1_11 <= reset ? 0 : _d__full_fsm___pip_5160_1_11;
_q__idx_fsm___pip_5160_1_12 <= reset ? 0 : _d__idx_fsm___pip_5160_1_12;
_q__full_fsm___pip_5160_1_12 <= reset ? 0 : _d__full_fsm___pip_5160_1_12;
_q__idx_fsm___pip_5160_1_13 <= reset ? 0 : _d__idx_fsm___pip_5160_1_13;
_q__full_fsm___pip_5160_1_13 <= reset ? 0 : _d__full_fsm___pip_5160_1_13;
_q__idx_fsm___pip_5160_1_14 <= reset ? 0 : _d__idx_fsm___pip_5160_1_14;
_q__full_fsm___pip_5160_1_14 <= reset ? 0 : _d__full_fsm___pip_5160_1_14;
_q__idx_fsm___pip_5160_1_15 <= reset ? 0 : _d__idx_fsm___pip_5160_1_15;
_q__full_fsm___pip_5160_1_15 <= reset ? 0 : _d__full_fsm___pip_5160_1_15;
_q__idx_fsm___pip_5160_1_16 <= reset ? 0 : _d__idx_fsm___pip_5160_1_16;
_q__full_fsm___pip_5160_1_16 <= reset ? 0 : _d__full_fsm___pip_5160_1_16;
_q__idx_fsm___pip_5160_1_17 <= reset ? 0 : _d__idx_fsm___pip_5160_1_17;
_q__full_fsm___pip_5160_1_17 <= reset ? 0 : _d__full_fsm___pip_5160_1_17;
_q__idx_fsm___pip_5160_1_18 <= reset ? 0 : _d__idx_fsm___pip_5160_1_18;
_q__full_fsm___pip_5160_1_18 <= reset ? 0 : _d__full_fsm___pip_5160_1_18;
_q__idx_fsm___pip_5160_1_19 <= reset ? 0 : _d__idx_fsm___pip_5160_1_19;
_q__full_fsm___pip_5160_1_19 <= reset ? 0 : _d__full_fsm___pip_5160_1_19;
_q__idx_fsm___pip_5160_1_20 <= reset ? 0 : _d__idx_fsm___pip_5160_1_20;
_q__full_fsm___pip_5160_1_20 <= reset ? 0 : _d__full_fsm___pip_5160_1_20;
_q__idx_fsm___pip_5160_1_21 <= reset ? 0 : _d__idx_fsm___pip_5160_1_21;
_q__full_fsm___pip_5160_1_21 <= reset ? 0 : _d__full_fsm___pip_5160_1_21;
_q__idx_fsm___pip_5160_1_22 <= reset ? 0 : _d__idx_fsm___pip_5160_1_22;
_q__full_fsm___pip_5160_1_22 <= reset ? 0 : _d__full_fsm___pip_5160_1_22;
_q__idx_fsm___pip_5160_1_23 <= reset ? 0 : _d__idx_fsm___pip_5160_1_23;
_q__full_fsm___pip_5160_1_23 <= reset ? 0 : _d__full_fsm___pip_5160_1_23;
_q__idx_fsm___pip_5160_1_24 <= reset ? 0 : _d__idx_fsm___pip_5160_1_24;
_q__full_fsm___pip_5160_1_24 <= reset ? 0 : _d__full_fsm___pip_5160_1_24;
_q__idx_fsm___pip_5160_1_25 <= reset ? 0 : _d__idx_fsm___pip_5160_1_25;
_q__full_fsm___pip_5160_1_25 <= reset ? 0 : _d__full_fsm___pip_5160_1_25;
_q__idx_fsm___pip_5160_1_26 <= reset ? 0 : _d__idx_fsm___pip_5160_1_26;
_q__full_fsm___pip_5160_1_26 <= reset ? 0 : _d__full_fsm___pip_5160_1_26;
_q__idx_fsm___pip_5160_1_27 <= reset ? 0 : _d__idx_fsm___pip_5160_1_27;
_q__full_fsm___pip_5160_1_27 <= reset ? 0 : _d__full_fsm___pip_5160_1_27;
_q__idx_fsm___pip_5160_1_28 <= reset ? 0 : _d__idx_fsm___pip_5160_1_28;
_q__full_fsm___pip_5160_1_28 <= reset ? 0 : _d__full_fsm___pip_5160_1_28;
_q__idx_fsm___pip_5160_1_29 <= reset ? 0 : _d__idx_fsm___pip_5160_1_29;
_q__full_fsm___pip_5160_1_29 <= reset ? 0 : _d__full_fsm___pip_5160_1_29;
_q__idx_fsm___pip_5160_1_30 <= reset ? 0 : _d__idx_fsm___pip_5160_1_30;
_q__full_fsm___pip_5160_1_30 <= reset ? 0 : _d__full_fsm___pip_5160_1_30;
_q__idx_fsm___pip_5160_1_31 <= reset ? 0 : _d__idx_fsm___pip_5160_1_31;
_q__full_fsm___pip_5160_1_31 <= reset ? 0 : _d__full_fsm___pip_5160_1_31;
_q__idx_fsm___pip_5160_1_32 <= reset ? 0 : _d__idx_fsm___pip_5160_1_32;
_q__full_fsm___pip_5160_1_32 <= reset ? 0 : _d__full_fsm___pip_5160_1_32;
_q__idx_fsm___pip_5160_1_33 <= reset ? 0 : _d__idx_fsm___pip_5160_1_33;
_q__full_fsm___pip_5160_1_33 <= reset ? 0 : _d__full_fsm___pip_5160_1_33;
_q__idx_fsm___pip_5160_1_34 <= reset ? 0 : _d__idx_fsm___pip_5160_1_34;
_q__full_fsm___pip_5160_1_34 <= reset ? 0 : _d__full_fsm___pip_5160_1_34;
_q__idx_fsm___pip_5160_1_35 <= reset ? 0 : _d__idx_fsm___pip_5160_1_35;
_q__full_fsm___pip_5160_1_35 <= reset ? 0 : _d__full_fsm___pip_5160_1_35;
_q__idx_fsm___pip_5160_1_36 <= reset ? 0 : _d__idx_fsm___pip_5160_1_36;
_q__full_fsm___pip_5160_1_36 <= reset ? 0 : _d__full_fsm___pip_5160_1_36;
_q__idx_fsm___pip_5160_1_37 <= reset ? 0 : _d__idx_fsm___pip_5160_1_37;
_q__full_fsm___pip_5160_1_37 <= reset ? 0 : _d__full_fsm___pip_5160_1_37;
_q__idx_fsm___pip_5160_1_38 <= reset ? 0 : _d__idx_fsm___pip_5160_1_38;
_q__full_fsm___pip_5160_1_38 <= reset ? 0 : _d__full_fsm___pip_5160_1_38;
_q__idx_fsm___pip_5160_1_39 <= reset ? 0 : _d__idx_fsm___pip_5160_1_39;
_q__full_fsm___pip_5160_1_39 <= reset ? 0 : _d__full_fsm___pip_5160_1_39;
_q__idx_fsm___pip_5160_1_40 <= reset ? 0 : _d__idx_fsm___pip_5160_1_40;
_q__full_fsm___pip_5160_1_40 <= reset ? 0 : _d__full_fsm___pip_5160_1_40;
_q__idx_fsm___pip_5160_1_41 <= reset ? 0 : _d__idx_fsm___pip_5160_1_41;
_q__full_fsm___pip_5160_1_41 <= reset ? 0 : _d__full_fsm___pip_5160_1_41;
_q__idx_fsm___pip_5160_1_42 <= reset ? 0 : _d__idx_fsm___pip_5160_1_42;
_q__full_fsm___pip_5160_1_42 <= reset ? 0 : _d__full_fsm___pip_5160_1_42;
_q__idx_fsm___pip_5160_1_43 <= reset ? 0 : _d__idx_fsm___pip_5160_1_43;
_q__full_fsm___pip_5160_1_43 <= reset ? 0 : _d__full_fsm___pip_5160_1_43;
_q__idx_fsm___pip_5160_1_44 <= reset ? 0 : _d__idx_fsm___pip_5160_1_44;
_q__full_fsm___pip_5160_1_44 <= reset ? 0 : _d__full_fsm___pip_5160_1_44;
_q__idx_fsm___pip_5160_1_45 <= reset ? 0 : _d__idx_fsm___pip_5160_1_45;
_q__full_fsm___pip_5160_1_45 <= reset ? 0 : _d__full_fsm___pip_5160_1_45;
_q__idx_fsm___pip_5160_1_46 <= reset ? 0 : _d__idx_fsm___pip_5160_1_46;
_q__full_fsm___pip_5160_1_46 <= reset ? 0 : _d__full_fsm___pip_5160_1_46;
_q__idx_fsm___pip_5160_1_47 <= reset ? 0 : _d__idx_fsm___pip_5160_1_47;
_q__full_fsm___pip_5160_1_47 <= reset ? 0 : _d__full_fsm___pip_5160_1_47;
_q__idx_fsm___pip_5160_1_48 <= reset ? 0 : _d__idx_fsm___pip_5160_1_48;
_q__full_fsm___pip_5160_1_48 <= reset ? 0 : _d__full_fsm___pip_5160_1_48;
_q__idx_fsm___pip_5160_1_49 <= reset ? 0 : _d__idx_fsm___pip_5160_1_49;
_q__full_fsm___pip_5160_1_49 <= reset ? 0 : _d__full_fsm___pip_5160_1_49;
_q__idx_fsm___pip_5160_1_50 <= reset ? 0 : _d__idx_fsm___pip_5160_1_50;
_q__full_fsm___pip_5160_1_50 <= reset ? 0 : _d__full_fsm___pip_5160_1_50;
_q__idx_fsm___pip_5160_1_51 <= reset ? 0 : _d__idx_fsm___pip_5160_1_51;
_q__full_fsm___pip_5160_1_51 <= reset ? 0 : _d__full_fsm___pip_5160_1_51;
_q__idx_fsm___pip_5160_1_52 <= reset ? 0 : _d__idx_fsm___pip_5160_1_52;
_q__full_fsm___pip_5160_1_52 <= reset ? 0 : _d__full_fsm___pip_5160_1_52;
_q__idx_fsm___pip_5160_1_53 <= reset ? 0 : _d__idx_fsm___pip_5160_1_53;
_q__full_fsm___pip_5160_1_53 <= reset ? 0 : _d__full_fsm___pip_5160_1_53;
_q__idx_fsm___pip_5160_1_54 <= reset ? 0 : _d__idx_fsm___pip_5160_1_54;
_q__full_fsm___pip_5160_1_54 <= reset ? 0 : _d__full_fsm___pip_5160_1_54;
_q__idx_fsm___pip_5160_1_55 <= reset ? 0 : _d__idx_fsm___pip_5160_1_55;
_q__full_fsm___pip_5160_1_55 <= reset ? 0 : _d__full_fsm___pip_5160_1_55;
_q__idx_fsm___pip_5160_1_56 <= reset ? 0 : _d__idx_fsm___pip_5160_1_56;
_q__full_fsm___pip_5160_1_56 <= reset ? 0 : _d__full_fsm___pip_5160_1_56;
_q__idx_fsm___pip_5160_1_57 <= reset ? 0 : _d__idx_fsm___pip_5160_1_57;
_q__full_fsm___pip_5160_1_57 <= reset ? 0 : _d__full_fsm___pip_5160_1_57;
_q__idx_fsm___pip_5160_1_58 <= reset ? 0 : _d__idx_fsm___pip_5160_1_58;
_q__full_fsm___pip_5160_1_58 <= reset ? 0 : _d__full_fsm___pip_5160_1_58;
_q__idx_fsm___pip_5160_1_59 <= reset ? 0 : _d__idx_fsm___pip_5160_1_59;
_q__full_fsm___pip_5160_1_59 <= reset ? 0 : _d__full_fsm___pip_5160_1_59;
_q__idx_fsm___pip_5160_1_60 <= reset ? 0 : _d__idx_fsm___pip_5160_1_60;
_q__full_fsm___pip_5160_1_60 <= reset ? 0 : _d__full_fsm___pip_5160_1_60;
_q__idx_fsm___pip_5160_1_61 <= reset ? 0 : _d__idx_fsm___pip_5160_1_61;
_q__full_fsm___pip_5160_1_61 <= reset ? 0 : _d__full_fsm___pip_5160_1_61;
_q__idx_fsm___pip_5160_1_62 <= reset ? 0 : _d__idx_fsm___pip_5160_1_62;
_q__full_fsm___pip_5160_1_62 <= reset ? 0 : _d__full_fsm___pip_5160_1_62;
_q__idx_fsm___pip_5160_1_63 <= reset ? 0 : _d__idx_fsm___pip_5160_1_63;
_q__full_fsm___pip_5160_1_63 <= reset ? 0 : _d__full_fsm___pip_5160_1_63;
_q__idx_fsm___pip_5160_1_64 <= reset ? 0 : _d__idx_fsm___pip_5160_1_64;
_q__full_fsm___pip_5160_1_64 <= reset ? 0 : _d__full_fsm___pip_5160_1_64;
_q__idx_fsm___pip_5160_1_65 <= reset ? 0 : _d__idx_fsm___pip_5160_1_65;
_q__full_fsm___pip_5160_1_65 <= reset ? 0 : _d__full_fsm___pip_5160_1_65;
_q__idx_fsm___pip_5160_1_66 <= reset ? 0 : _d__idx_fsm___pip_5160_1_66;
_q__full_fsm___pip_5160_1_66 <= reset ? 0 : _d__full_fsm___pip_5160_1_66;
_q__idx_fsm___pip_5160_1_67 <= reset ? 0 : _d__idx_fsm___pip_5160_1_67;
_q__full_fsm___pip_5160_1_67 <= reset ? 0 : _d__full_fsm___pip_5160_1_67;
_q__idx_fsm___pip_5160_1_68 <= reset ? 0 : _d__idx_fsm___pip_5160_1_68;
_q__full_fsm___pip_5160_1_68 <= reset ? 0 : _d__full_fsm___pip_5160_1_68;
_q__idx_fsm___pip_5160_1_69 <= reset ? 0 : _d__idx_fsm___pip_5160_1_69;
_q__full_fsm___pip_5160_1_69 <= reset ? 0 : _d__full_fsm___pip_5160_1_69;
_q__idx_fsm___pip_5160_1_70 <= reset ? 0 : _d__idx_fsm___pip_5160_1_70;
_q__full_fsm___pip_5160_1_70 <= reset ? 0 : _d__full_fsm___pip_5160_1_70;
_q__idx_fsm___pip_5160_1_71 <= reset ? 0 : _d__idx_fsm___pip_5160_1_71;
_q__full_fsm___pip_5160_1_71 <= reset ? 0 : _d__full_fsm___pip_5160_1_71;
_q__idx_fsm___pip_5160_1_72 <= reset ? 0 : _d__idx_fsm___pip_5160_1_72;
_q__full_fsm___pip_5160_1_72 <= reset ? 0 : _d__full_fsm___pip_5160_1_72;
_q__idx_fsm___pip_5160_1_73 <= reset ? 0 : _d__idx_fsm___pip_5160_1_73;
_q__full_fsm___pip_5160_1_73 <= reset ? 0 : _d__full_fsm___pip_5160_1_73;
_q__idx_fsm___pip_5160_1_74 <= reset ? 0 : _d__idx_fsm___pip_5160_1_74;
_q__full_fsm___pip_5160_1_74 <= reset ? 0 : _d__full_fsm___pip_5160_1_74;
_q__idx_fsm___pip_5160_1_75 <= reset ? 0 : _d__idx_fsm___pip_5160_1_75;
_q__full_fsm___pip_5160_1_75 <= reset ? 0 : _d__full_fsm___pip_5160_1_75;
_q__idx_fsm___pip_5160_1_76 <= reset ? 0 : _d__idx_fsm___pip_5160_1_76;
_q__full_fsm___pip_5160_1_76 <= reset ? 0 : _d__full_fsm___pip_5160_1_76;
_q__idx_fsm___pip_5160_1_77 <= reset ? 0 : _d__idx_fsm___pip_5160_1_77;
_q__full_fsm___pip_5160_1_77 <= reset ? 0 : _d__full_fsm___pip_5160_1_77;
_q__idx_fsm___pip_5160_1_78 <= reset ? 0 : _d__idx_fsm___pip_5160_1_78;
_q__full_fsm___pip_5160_1_78 <= reset ? 0 : _d__full_fsm___pip_5160_1_78;
_q__idx_fsm___pip_5160_1_79 <= reset ? 0 : _d__idx_fsm___pip_5160_1_79;
_q__full_fsm___pip_5160_1_79 <= reset ? 0 : _d__full_fsm___pip_5160_1_79;
_q__idx_fsm___pip_5160_1_80 <= reset ? 0 : _d__idx_fsm___pip_5160_1_80;
_q__full_fsm___pip_5160_1_80 <= reset ? 0 : _d__full_fsm___pip_5160_1_80;
_q__idx_fsm___pip_5160_1_81 <= reset ? 0 : _d__idx_fsm___pip_5160_1_81;
_q__full_fsm___pip_5160_1_81 <= reset ? 0 : _d__full_fsm___pip_5160_1_81;
_q__idx_fsm___pip_5160_1_82 <= reset ? 0 : _d__idx_fsm___pip_5160_1_82;
_q__full_fsm___pip_5160_1_82 <= reset ? 0 : _d__full_fsm___pip_5160_1_82;
_q__idx_fsm___pip_5160_1_83 <= reset ? 0 : _d__idx_fsm___pip_5160_1_83;
_q__full_fsm___pip_5160_1_83 <= reset ? 0 : _d__full_fsm___pip_5160_1_83;
_q__idx_fsm___pip_5160_1_84 <= reset ? 0 : _d__idx_fsm___pip_5160_1_84;
_q__full_fsm___pip_5160_1_84 <= reset ? 0 : _d__full_fsm___pip_5160_1_84;
_q__idx_fsm___pip_5160_1_85 <= reset ? 0 : _d__idx_fsm___pip_5160_1_85;
_q__full_fsm___pip_5160_1_85 <= reset ? 0 : _d__full_fsm___pip_5160_1_85;
_q__idx_fsm___pip_5160_1_86 <= reset ? 0 : _d__idx_fsm___pip_5160_1_86;
_q__full_fsm___pip_5160_1_86 <= reset ? 0 : _d__full_fsm___pip_5160_1_86;
_q__idx_fsm___pip_5160_1_87 <= reset ? 0 : _d__idx_fsm___pip_5160_1_87;
_q__full_fsm___pip_5160_1_87 <= reset ? 0 : _d__full_fsm___pip_5160_1_87;
_q__idx_fsm___pip_5160_1_88 <= reset ? 0 : _d__idx_fsm___pip_5160_1_88;
_q__full_fsm___pip_5160_1_88 <= reset ? 0 : _d__full_fsm___pip_5160_1_88;
_q__idx_fsm___pip_5160_1_89 <= reset ? 0 : _d__idx_fsm___pip_5160_1_89;
_q__full_fsm___pip_5160_1_89 <= reset ? 0 : _d__full_fsm___pip_5160_1_89;
_q__idx_fsm___pip_5160_1_90 <= reset ? 0 : _d__idx_fsm___pip_5160_1_90;
_q__full_fsm___pip_5160_1_90 <= reset ? 0 : _d__full_fsm___pip_5160_1_90;
_q__idx_fsm___pip_5160_1_91 <= reset ? 0 : _d__idx_fsm___pip_5160_1_91;
_q__full_fsm___pip_5160_1_91 <= reset ? 0 : _d__full_fsm___pip_5160_1_91;
_q__idx_fsm___pip_5160_1_92 <= reset ? 0 : _d__idx_fsm___pip_5160_1_92;
_q__full_fsm___pip_5160_1_92 <= reset ? 0 : _d__full_fsm___pip_5160_1_92;
_q__idx_fsm___pip_5160_1_93 <= reset ? 0 : _d__idx_fsm___pip_5160_1_93;
_q__full_fsm___pip_5160_1_93 <= reset ? 0 : _d__full_fsm___pip_5160_1_93;
_q__idx_fsm___pip_5160_1_94 <= reset ? 0 : _d__idx_fsm___pip_5160_1_94;
_q__full_fsm___pip_5160_1_94 <= reset ? 0 : _d__full_fsm___pip_5160_1_94;
_q__idx_fsm___pip_5160_1_95 <= reset ? 0 : _d__idx_fsm___pip_5160_1_95;
_q__full_fsm___pip_5160_1_95 <= reset ? 0 : _d__full_fsm___pip_5160_1_95;
_q__idx_fsm___pip_5160_1_96 <= reset ? 0 : _d__idx_fsm___pip_5160_1_96;
_q__full_fsm___pip_5160_1_96 <= reset ? 0 : _d__full_fsm___pip_5160_1_96;
_q__idx_fsm___pip_5160_1_97 <= reset ? 0 : _d__idx_fsm___pip_5160_1_97;
_q__full_fsm___pip_5160_1_97 <= reset ? 0 : _d__full_fsm___pip_5160_1_97;
_q__idx_fsm___pip_5160_1_98 <= reset ? 0 : _d__idx_fsm___pip_5160_1_98;
_q__full_fsm___pip_5160_1_98 <= reset ? 0 : _d__full_fsm___pip_5160_1_98;
_q__idx_fsm___pip_5160_1_99 <= reset ? 0 : _d__idx_fsm___pip_5160_1_99;
_q__full_fsm___pip_5160_1_99 <= reset ? 0 : _d__full_fsm___pip_5160_1_99;
_q__idx_fsm___pip_5160_1_100 <= reset ? 0 : _d__idx_fsm___pip_5160_1_100;
_q__full_fsm___pip_5160_1_100 <= reset ? 0 : _d__full_fsm___pip_5160_1_100;
_q__idx_fsm___pip_5160_1_101 <= reset ? 0 : _d__idx_fsm___pip_5160_1_101;
_q__full_fsm___pip_5160_1_101 <= reset ? 0 : _d__full_fsm___pip_5160_1_101;
_q__idx_fsm___pip_5160_1_102 <= reset ? 0 : _d__idx_fsm___pip_5160_1_102;
_q__full_fsm___pip_5160_1_102 <= reset ? 0 : _d__full_fsm___pip_5160_1_102;
_q__idx_fsm___pip_5160_1_103 <= reset ? 0 : _d__idx_fsm___pip_5160_1_103;
_q__full_fsm___pip_5160_1_103 <= reset ? 0 : _d__full_fsm___pip_5160_1_103;
_q__idx_fsm___pip_5160_1_104 <= reset ? 0 : _d__idx_fsm___pip_5160_1_104;
_q__full_fsm___pip_5160_1_104 <= reset ? 0 : _d__full_fsm___pip_5160_1_104;
_q__idx_fsm___pip_5160_1_105 <= reset ? 0 : _d__idx_fsm___pip_5160_1_105;
_q__full_fsm___pip_5160_1_105 <= reset ? 0 : _d__full_fsm___pip_5160_1_105;
_q__idx_fsm___pip_5160_1_106 <= reset ? 0 : _d__idx_fsm___pip_5160_1_106;
_q__full_fsm___pip_5160_1_106 <= reset ? 0 : _d__full_fsm___pip_5160_1_106;
_q__idx_fsm___pip_5160_1_107 <= reset ? 0 : _d__idx_fsm___pip_5160_1_107;
_q__full_fsm___pip_5160_1_107 <= reset ? 0 : _d__full_fsm___pip_5160_1_107;
_q__idx_fsm___pip_5160_1_108 <= reset ? 0 : _d__idx_fsm___pip_5160_1_108;
_q__full_fsm___pip_5160_1_108 <= reset ? 0 : _d__full_fsm___pip_5160_1_108;
_q__idx_fsm___pip_5160_1_109 <= reset ? 0 : _d__idx_fsm___pip_5160_1_109;
_q__full_fsm___pip_5160_1_109 <= reset ? 0 : _d__full_fsm___pip_5160_1_109;
_q__idx_fsm___pip_5160_1_110 <= reset ? 0 : _d__idx_fsm___pip_5160_1_110;
_q__full_fsm___pip_5160_1_110 <= reset ? 0 : _d__full_fsm___pip_5160_1_110;
_q__idx_fsm___pip_5160_1_111 <= reset ? 0 : _d__idx_fsm___pip_5160_1_111;
_q__full_fsm___pip_5160_1_111 <= reset ? 0 : _d__full_fsm___pip_5160_1_111;
_q__idx_fsm___pip_5160_1_112 <= reset ? 0 : _d__idx_fsm___pip_5160_1_112;
_q__full_fsm___pip_5160_1_112 <= reset ? 0 : _d__full_fsm___pip_5160_1_112;
_q__idx_fsm___pip_5160_1_113 <= reset ? 0 : _d__idx_fsm___pip_5160_1_113;
_q__full_fsm___pip_5160_1_113 <= reset ? 0 : _d__full_fsm___pip_5160_1_113;
_q__idx_fsm___pip_5160_1_114 <= reset ? 0 : _d__idx_fsm___pip_5160_1_114;
_q__full_fsm___pip_5160_1_114 <= reset ? 0 : _d__full_fsm___pip_5160_1_114;
_q__idx_fsm___pip_5160_1_115 <= reset ? 0 : _d__idx_fsm___pip_5160_1_115;
_q__full_fsm___pip_5160_1_115 <= reset ? 0 : _d__full_fsm___pip_5160_1_115;
_q__idx_fsm___pip_5160_1_116 <= reset ? 0 : _d__idx_fsm___pip_5160_1_116;
_q__full_fsm___pip_5160_1_116 <= reset ? 0 : _d__full_fsm___pip_5160_1_116;
_q__idx_fsm___pip_5160_1_117 <= reset ? 0 : _d__idx_fsm___pip_5160_1_117;
_q__full_fsm___pip_5160_1_117 <= reset ? 0 : _d__full_fsm___pip_5160_1_117;
_q__idx_fsm___pip_5160_1_118 <= reset ? 0 : _d__idx_fsm___pip_5160_1_118;
_q__full_fsm___pip_5160_1_118 <= reset ? 0 : _d__full_fsm___pip_5160_1_118;
_q__idx_fsm___pip_5160_1_119 <= reset ? 0 : _d__idx_fsm___pip_5160_1_119;
_q__full_fsm___pip_5160_1_119 <= reset ? 0 : _d__full_fsm___pip_5160_1_119;
_q__idx_fsm___pip_5160_1_120 <= reset ? 0 : _d__idx_fsm___pip_5160_1_120;
_q__full_fsm___pip_5160_1_120 <= reset ? 0 : _d__full_fsm___pip_5160_1_120;
_q__idx_fsm___pip_5160_1_121 <= reset ? 0 : _d__idx_fsm___pip_5160_1_121;
_q__full_fsm___pip_5160_1_121 <= reset ? 0 : _d__full_fsm___pip_5160_1_121;
_q__idx_fsm___pip_5160_1_122 <= reset ? 0 : _d__idx_fsm___pip_5160_1_122;
_q__full_fsm___pip_5160_1_122 <= reset ? 0 : _d__full_fsm___pip_5160_1_122;
_q__idx_fsm___pip_5160_1_123 <= reset ? 0 : _d__idx_fsm___pip_5160_1_123;
_q__full_fsm___pip_5160_1_123 <= reset ? 0 : _d__full_fsm___pip_5160_1_123;
_q__idx_fsm___pip_5160_1_124 <= reset ? 0 : _d__idx_fsm___pip_5160_1_124;
_q__full_fsm___pip_5160_1_124 <= reset ? 0 : _d__full_fsm___pip_5160_1_124;
_q__idx_fsm___pip_5160_1_125 <= reset ? 0 : _d__idx_fsm___pip_5160_1_125;
_q__full_fsm___pip_5160_1_125 <= reset ? 0 : _d__full_fsm___pip_5160_1_125;
_q__idx_fsm___pip_5160_1_126 <= reset ? 0 : _d__idx_fsm___pip_5160_1_126;
_q__full_fsm___pip_5160_1_126 <= reset ? 0 : _d__full_fsm___pip_5160_1_126;
_q__idx_fsm___pip_5160_1_127 <= reset ? 0 : _d__idx_fsm___pip_5160_1_127;
_q__full_fsm___pip_5160_1_127 <= reset ? 0 : _d__full_fsm___pip_5160_1_127;
_q__idx_fsm___pip_5160_1_128 <= reset ? 0 : _d__idx_fsm___pip_5160_1_128;
_q__full_fsm___pip_5160_1_128 <= reset ? 0 : _d__full_fsm___pip_5160_1_128;
_q__idx_fsm___pip_5160_1_129 <= reset ? 0 : _d__idx_fsm___pip_5160_1_129;
_q__full_fsm___pip_5160_1_129 <= reset ? 0 : _d__full_fsm___pip_5160_1_129;
_q__idx_fsm___pip_5160_1_130 <= reset ? 0 : _d__idx_fsm___pip_5160_1_130;
_q__full_fsm___pip_5160_1_130 <= reset ? 0 : _d__full_fsm___pip_5160_1_130;
_q__idx_fsm___pip_5160_1_131 <= reset ? 0 : _d__idx_fsm___pip_5160_1_131;
_q__full_fsm___pip_5160_1_131 <= reset ? 0 : _d__full_fsm___pip_5160_1_131;
_q__idx_fsm___pip_5160_1_132 <= reset ? 0 : _d__idx_fsm___pip_5160_1_132;
_q__full_fsm___pip_5160_1_132 <= reset ? 0 : _d__full_fsm___pip_5160_1_132;
_q__idx_fsm___pip_5160_1_133 <= reset ? 0 : _d__idx_fsm___pip_5160_1_133;
_q__full_fsm___pip_5160_1_133 <= reset ? 0 : _d__full_fsm___pip_5160_1_133;
_q__idx_fsm___pip_5160_1_134 <= reset ? 0 : _d__idx_fsm___pip_5160_1_134;
_q__full_fsm___pip_5160_1_134 <= reset ? 0 : _d__full_fsm___pip_5160_1_134;
_q__idx_fsm___pip_5160_1_135 <= reset ? 0 : _d__idx_fsm___pip_5160_1_135;
_q__full_fsm___pip_5160_1_135 <= reset ? 0 : _d__full_fsm___pip_5160_1_135;
_q__idx_fsm___pip_5160_1_136 <= reset ? 0 : _d__idx_fsm___pip_5160_1_136;
_q__full_fsm___pip_5160_1_136 <= reset ? 0 : _d__full_fsm___pip_5160_1_136;
end

endmodule


projf-explore/lib/memory/rom_async.sv
projf-explore/lib/memory/bram_sdp.sv